module interrupt_priority_resolve (
	clk,
	n_rst,
	interrupt_priorities,
	pending_interrupts,
	active_interrupt,
	active_interrupt_ID,
	interrupt_processing
);
	parameter N_INTERRUPTS = 32;
	input wire clk;
	input wire n_rst;
	input wire [(N_INTERRUPTS * 32) - 1:0] interrupt_priorities;
	input wire [N_INTERRUPTS - 1:0] pending_interrupts;
	output wire [N_INTERRUPTS - 1:0] active_interrupt;
	output wire [31:0] active_interrupt_ID;
	output wire interrupt_processing;
	wire [(N_INTERRUPTS * 32) - 1:0] max_ids;
	wire [(N_INTERRUPTS * 32) - 1:0] max_priorities;
	wire [(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? (((($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) - ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS)) + 1) * 32) + ((($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) * 32) - 1) : (((($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1))) + 1) * 32) + ((($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) * 32) - 1)):(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) * 32 : ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) * 32)] ids;
	wire [(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? (((($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) - ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS)) + 1) * 32) + ((($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) * 32) - 1) : (((($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1))) + 1) * 32) + ((($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) * 32) - 1)):(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) * 32 : ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) * 32)] priorities;
	wire interrupt_process;
	reg interrupt_process_prev;
	assign active_interrupt_ID = (ids[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? ($clog2(N_INTERRUPTS) >= 0 ? $clog2(N_INTERRUPTS) : $clog2(N_INTERRUPTS) - $clog2(N_INTERRUPTS)) * N_INTERRUPTS : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - ((($clog2(N_INTERRUPTS) >= 0 ? $clog2(N_INTERRUPTS) : $clog2(N_INTERRUPTS) - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32] == 0 ? {32 {1'sb0}} : ids[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? ($clog2(N_INTERRUPTS) >= 0 ? $clog2(N_INTERRUPTS) : $clog2(N_INTERRUPTS) - $clog2(N_INTERRUPTS)) * N_INTERRUPTS : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - ((($clog2(N_INTERRUPTS) >= 0 ? $clog2(N_INTERRUPTS) : $clog2(N_INTERRUPTS) - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32]);
	assign active_interrupt = (ids[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? ($clog2(N_INTERRUPTS) >= 0 ? $clog2(N_INTERRUPTS) : $clog2(N_INTERRUPTS) - $clog2(N_INTERRUPTS)) * N_INTERRUPTS : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - ((($clog2(N_INTERRUPTS) >= 0 ? $clog2(N_INTERRUPTS) : $clog2(N_INTERRUPTS) - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32] == 0 ? {N_INTERRUPTS {1'sb0}} : 'b1 << (ids[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? ($clog2(N_INTERRUPTS) >= 0 ? $clog2(N_INTERRUPTS) : $clog2(N_INTERRUPTS) - $clog2(N_INTERRUPTS)) * N_INTERRUPTS : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - ((($clog2(N_INTERRUPTS) >= 0 ? $clog2(N_INTERRUPTS) : $clog2(N_INTERRUPTS) - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32] - 1));
	assign interrupt_process = pending_interrupts != {N_INTERRUPTS {1'sb0}};
	assign interrupt_processing = interrupt_process & ~interrupt_process_prev;
	always @(posedge clk or negedge n_rst)
		if (!n_rst)
			interrupt_process_prev <= 1'b0;
		else
			interrupt_process_prev <= interrupt_process;
	genvar i;
	genvar j;
	generate
		for (i = 0; i <= $clog2(N_INTERRUPTS); i = i + 1) for (j = 0; j < (2 ** ($clog2(N_INTERRUPTS) - i)); j = j + 1) if (i == 0) begin
			assign ids[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? (($clog2(N_INTERRUPTS) >= 0 ? i : $clog2(N_INTERRUPTS) - i) * N_INTERRUPTS) + j : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - (((($clog2(N_INTERRUPTS) >= 0 ? i : $clog2(N_INTERRUPTS) - i) * N_INTERRUPTS) + j) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32] = (pending_interrupts[j] ? j + 1 : 0);
			assign priorities[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? (($clog2(N_INTERRUPTS) >= 0 ? i : $clog2(N_INTERRUPTS) - i) * N_INTERRUPTS) + j : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - (((($clog2(N_INTERRUPTS) >= 0 ? i : $clog2(N_INTERRUPTS) - i) * N_INTERRUPTS) + j) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32] = (pending_interrupts[j] ? interrupt_priorities[j * 32+:32] : 0);
		end
		else begin
			assign ids[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? (($clog2(N_INTERRUPTS) >= 0 ? i : $clog2(N_INTERRUPTS) - i) * N_INTERRUPTS) + j : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - (((($clog2(N_INTERRUPTS) >= 0 ? i : $clog2(N_INTERRUPTS) - i) * N_INTERRUPTS) + j) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32] = (priorities[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? (($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + (2 * j) : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - (((($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + (2 * j)) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32] >= priorities[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? (($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + ((2 * j) + 1) : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - (((($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + ((2 * j) + 1)) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32] ? ids[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? (($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + (2 * j) : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - (((($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + (2 * j)) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32] : ids[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? (($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + ((2 * j) + 1) : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - (((($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + ((2 * j) + 1)) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32]);
			assign priorities[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? (($clog2(N_INTERRUPTS) >= 0 ? i : $clog2(N_INTERRUPTS) - i) * N_INTERRUPTS) + j : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - (((($clog2(N_INTERRUPTS) >= 0 ? i : $clog2(N_INTERRUPTS) - i) * N_INTERRUPTS) + j) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32] = (priorities[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? (($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + (2 * j) : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - (((($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + (2 * j)) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32] >= priorities[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? (($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + ((2 * j) + 1) : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - (((($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + ((2 * j) + 1)) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32] ? priorities[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? (($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + (2 * j) : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - (((($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + (2 * j)) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32] : priorities[(($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)) >= ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) ? (($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + ((2 * j) + 1) : ($clog2(N_INTERRUPTS) >= 0 ? 0 : $clog2(N_INTERRUPTS) * N_INTERRUPTS) - (((($clog2(N_INTERRUPTS) >= 0 ? i - 1 : $clog2(N_INTERRUPTS) - (i - 1)) * N_INTERRUPTS) + ((2 * j) + 1)) - ($clog2(N_INTERRUPTS) >= 0 ? (($clog2(N_INTERRUPTS) + 1) * N_INTERRUPTS) - 1 : ((1 - $clog2(N_INTERRUPTS)) * N_INTERRUPTS) + (($clog2(N_INTERRUPTS) * N_INTERRUPTS) - 1)))) * 32+:32]);
		end
	endgenerate
endmodule

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_level_bASIC
  CLASS BLOCK ;
  FOREIGN top_level_bASIC ;
  ORIGIN 0.000 0.000 ;
  SIZE 2700.000 BY 3300.000 ;
  PIN MISO_bi
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2616.110 0.000 2616.390 4.000 ;
    END
  END MISO_bi
  PIN MISO_output_en_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.610 0.000 2627.890 4.000 ;
    END
  END MISO_output_en_low
  PIN MOSI_bi
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END MOSI_bi
  PIN MOSI_output_en_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.650 0.000 2638.930 4.000 ;
    END
  END MOSI_output_en_low
  PIN SCK_bi
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 3296.000 96.510 3300.000 ;
    END
  END SCK_bi
  PIN SCK_output_en_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 274.760 2700.000 275.360 ;
    END
  END SCK_output_en_low
  PIN SCL_bi
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 3296.000 289.250 3300.000 ;
    END
  END SCL_bi
  PIN SCL_output_en_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END SCL_output_en_low
  PIN SDA_bi
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 3296.000 481.990 3300.000 ;
    END
  END SDA_bi
  PIN SDA_output_en_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 824.200 2700.000 824.800 ;
    END
  END SDA_output_en_low
  PIN SS_bi
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 3296.000 674.730 3300.000 ;
    END
  END SS_bi
  PIN SS_output_en_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2649.690 0.000 2649.970 4.000 ;
    END
  END SS_output_en_low
  PIN asyncrst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.650 3296.000 867.930 3300.000 ;
    END
  END asyncrst_n
  PIN clk_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END clk_sel
  PIN gpio_bidir_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.130 3296.000 1253.410 3300.000 ;
    END
  END gpio_bidir_io[0]
  PIN gpio_bidir_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.070 3296.000 1639.350 3300.000 ;
    END
  END gpio_bidir_io[1]
  PIN gpio_bidir_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2249.480 4.000 2250.080 ;
    END
  END gpio_bidir_io[2]
  PIN gpio_bidir_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1831.810 3296.000 1832.090 3300.000 ;
    END
  END gpio_bidir_io[3]
  PIN gpio_bidir_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2217.750 3296.000 2218.030 3300.000 ;
    END
  END gpio_bidir_io[4]
  PIN gpio_bidir_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2474.560 2700.000 2475.160 ;
    END
  END gpio_bidir_io[5]
  PIN gpio_bidir_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3024.680 2700.000 3025.280 ;
    END
  END gpio_bidir_io[6]
  PIN gpio_bidir_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.230 3296.000 2603.510 3300.000 ;
    END
  END gpio_bidir_io[7]
  PIN gpio_output_en_low[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.330 3296.000 1446.610 3300.000 ;
    END
  END gpio_output_en_low[0]
  PIN gpio_output_en_low[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1649.040 4.000 1649.640 ;
    END
  END gpio_output_en_low[1]
  PIN gpio_output_en_low[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2683.270 0.000 2683.550 4.000 ;
    END
  END gpio_output_en_low[2]
  PIN gpio_output_en_low[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2024.550 3296.000 2024.830 3300.000 ;
    END
  END gpio_output_en_low[3]
  PIN gpio_output_en_low[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2410.490 3296.000 2410.770 3300.000 ;
    END
  END gpio_output_en_low[4]
  PIN gpio_output_en_low[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2849.240 4.000 2849.840 ;
    END
  END gpio_output_en_low[5]
  PIN gpio_output_en_low[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2694.310 0.000 2694.590 4.000 ;
    END
  END gpio_output_en_low[6]
  PIN gpio_output_en_low[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3149.120 4.000 3149.720 ;
    END
  END gpio_output_en_low[7]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1924.440 2700.000 1925.040 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1949.600 4.000 1950.200 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2549.360 4.000 2549.960 ;
    END
  END irq[2]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 0.000 1188.550 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2303.770 0.000 2304.050 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2315.270 0.000 2315.550 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2326.310 0.000 2326.590 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.350 0.000 2337.630 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2348.390 0.000 2348.670 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2359.890 0.000 2360.170 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2370.930 0.000 2371.210 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2381.970 0.000 2382.250 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2393.010 0.000 2393.290 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2404.510 0.000 2404.790 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.590 0.000 1299.870 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2415.550 0.000 2415.830 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2426.590 0.000 2426.870 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.630 0.000 2437.910 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.130 0.000 2449.410 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2460.170 0.000 2460.450 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2471.210 0.000 2471.490 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2482.250 0.000 2482.530 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2493.750 0.000 2494.030 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2504.790 0.000 2505.070 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2515.830 0.000 2516.110 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 0.000 1310.910 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.870 0.000 2527.150 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.370 0.000 2538.650 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2549.410 0.000 2549.690 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2560.450 0.000 2560.730 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.490 0.000 2571.770 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2582.990 0.000 2583.270 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2594.030 0.000 2594.310 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2605.070 0.000 2605.350 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.130 0.000 1322.410 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.170 0.000 1333.450 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.210 0.000 1344.490 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 0.000 1355.990 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.750 0.000 1367.030 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.790 0.000 1378.070 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.830 0.000 1389.110 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.330 0.000 1400.610 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.310 0.000 1199.590 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1411.370 0.000 1411.650 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.410 0.000 1422.690 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.450 0.000 1433.730 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.950 0.000 1445.230 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.990 0.000 1456.270 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.030 0.000 1467.310 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.070 0.000 1478.350 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.570 0.000 1489.850 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.610 0.000 1500.890 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.650 0.000 1511.930 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.350 0.000 1210.630 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.690 0.000 1522.970 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.190 0.000 1534.470 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.230 0.000 1545.510 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1556.270 0.000 1556.550 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.310 0.000 1567.590 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.810 0.000 1579.090 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.850 0.000 1590.130 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.890 0.000 1601.170 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.930 0.000 1612.210 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1623.430 0.000 1623.710 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.390 0.000 1221.670 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.470 0.000 1634.750 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.510 0.000 1645.790 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.550 0.000 1656.830 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.050 0.000 1668.330 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.090 0.000 1679.370 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.130 0.000 1690.410 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1701.170 0.000 1701.450 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.670 0.000 1712.950 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1723.710 0.000 1723.990 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.750 0.000 1735.030 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.890 0.000 1233.170 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.790 0.000 1746.070 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1757.290 0.000 1757.570 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.330 0.000 1768.610 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1779.370 0.000 1779.650 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.410 0.000 1790.690 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1801.910 0.000 1802.190 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.950 0.000 1813.230 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.990 0.000 1824.270 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.490 0.000 1835.770 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.530 0.000 1846.810 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.930 0.000 1244.210 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.570 0.000 1857.850 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.610 0.000 1868.890 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1880.110 0.000 1880.390 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1891.150 0.000 1891.430 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1902.190 0.000 1902.470 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1913.230 0.000 1913.510 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1924.730 0.000 1925.010 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.770 0.000 1936.050 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1946.810 0.000 1947.090 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1957.850 0.000 1958.130 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1254.970 0.000 1255.250 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1969.350 0.000 1969.630 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.390 0.000 1980.670 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1991.430 0.000 1991.710 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2002.470 0.000 2002.750 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2013.970 0.000 2014.250 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.010 0.000 2025.290 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.050 0.000 2036.330 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.090 0.000 2047.370 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2058.590 0.000 2058.870 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2069.630 0.000 2069.910 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.010 0.000 1266.290 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.670 0.000 2080.950 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2091.710 0.000 2091.990 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2103.210 0.000 2103.490 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2114.250 0.000 2114.530 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.290 0.000 2125.570 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.330 0.000 2136.610 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.830 0.000 2148.110 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2158.870 0.000 2159.150 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2169.910 0.000 2170.190 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.950 0.000 2181.230 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.510 0.000 1277.790 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2192.450 0.000 2192.730 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2203.490 0.000 2203.770 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2214.530 0.000 2214.810 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2225.570 0.000 2225.850 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2237.070 0.000 2237.350 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.110 0.000 2248.390 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2259.150 0.000 2259.430 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2270.650 0.000 2270.930 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2281.690 0.000 2281.970 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.730 0.000 2293.010 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.550 0.000 1288.830 4.000 ;
    END
  END la_data_out[9]
  PIN pwm_w_data_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1049.280 4.000 1049.880 ;
    END
  END pwm_w_data_0
  PIN timer_bidir_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2660.730 0.000 2661.010 4.000 ;
    END
  END timer_bidir_0
  PIN timer_output_en_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2672.230 0.000 2672.510 4.000 ;
    END
  END timer_output_en_low
  PIN uart_debug_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1374.320 2700.000 1374.920 ;
    END
  END uart_debug_rx
  PIN uart_debug_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.160 4.000 1349.760 ;
    END
  END uart_debug_tx
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.390 3296.000 1060.670 3300.000 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.250 0.000 619.530 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 0.000 652.650 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 0.000 719.810 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.110 0.000 753.390 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 0.000 786.510 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 0.000 820.090 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.970 0.000 887.250 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 0.000 920.830 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.670 0.000 953.950 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 0.000 987.530 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.410 0.000 1054.690 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.530 0.000 1087.810 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.110 0.000 1121.390 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.690 0.000 1154.970 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 0.000 563.410 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 0.000 596.990 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 0.000 630.570 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 0.000 697.270 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 0.000 730.850 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.150 0.000 764.430 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 0.000 798.010 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.430 0.000 864.710 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.010 0.000 898.290 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.590 0.000 931.870 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.170 0.000 965.450 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 0.000 998.570 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.870 0.000 1032.150 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.450 0.000 1065.730 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.030 0.000 1099.310 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.150 0.000 1132.430 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 0.000 1166.010 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.750 0.000 608.030 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 0.000 641.610 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 0.000 741.890 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 0.000 775.470 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.770 0.000 809.050 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 0.000 842.630 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.470 0.000 875.750 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.050 0.000 909.330 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.630 0.000 942.910 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.210 0.000 976.490 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.790 0.000 1010.070 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.910 0.000 1043.190 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.490 0.000 1076.770 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.070 0.000 1110.350 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.650 0.000 1143.930 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.770 0.000 1177.050 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 3171.070 2633.840 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 3171.070 2480.240 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 3171.070 2326.640 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 3171.070 2173.040 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 3171.070 2019.440 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 2657.930 2633.840 2738.410 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 2657.930 2480.240 2738.410 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 2657.930 2326.640 2738.410 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 2657.930 2173.040 2738.410 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 2657.930 2019.440 2738.410 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 2144.790 2633.840 2225.270 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 2144.790 2480.240 2225.270 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 2144.790 2326.640 2225.270 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 2144.790 2173.040 2225.270 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 2144.790 2019.440 2225.270 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 1631.650 2633.840 1712.130 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 1631.650 2480.240 1712.130 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 1631.650 2326.640 1712.130 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 1631.650 2173.040 1712.130 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 1631.650 2019.440 1712.130 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 1118.510 2633.840 1198.990 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 1118.510 2480.240 1198.990 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 1118.510 2326.640 1198.990 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 1118.510 2173.040 1198.990 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 1118.510 2019.440 1198.990 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 605.370 2633.840 685.850 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 605.370 2480.240 685.850 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 605.370 2326.640 685.850 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 605.370 2173.040 685.850 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 605.370 2019.440 685.850 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 172.710 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 172.710 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 172.710 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 172.710 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 172.710 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 3171.070 2557.040 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 3171.070 2403.440 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 3171.070 2249.840 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 3171.070 2096.240 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 2657.930 2557.040 2738.410 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 2657.930 2403.440 2738.410 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 2657.930 2249.840 2738.410 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 2657.930 2096.240 2738.410 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 2144.790 2557.040 2225.270 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 2144.790 2403.440 2225.270 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 2144.790 2249.840 2225.270 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 2144.790 2096.240 2225.270 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 1631.650 2557.040 1712.130 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 1631.650 2403.440 1712.130 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 1631.650 2249.840 1712.130 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 1631.650 2096.240 1712.130 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 1118.510 2557.040 1198.990 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 1118.510 2403.440 1198.990 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 1118.510 2249.840 1198.990 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 1118.510 2096.240 1198.990 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 605.370 2557.040 685.850 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 605.370 2403.440 685.850 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 605.370 2249.840 685.850 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 605.370 2096.240 685.850 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 172.710 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 172.710 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 172.710 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 172.710 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2635.540 3171.310 2637.140 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2481.940 3171.310 2483.540 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2328.340 3171.310 2329.940 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2174.740 3171.310 2176.340 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.140 3171.310 2022.740 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1867.540 10.880 1869.140 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1713.940 10.880 1715.540 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1560.340 10.880 1561.940 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1406.740 10.880 1408.340 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1253.140 10.880 1254.740 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1099.540 10.880 1101.140 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 945.940 10.880 947.540 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.340 10.880 793.940 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2635.540 2658.170 2637.140 2738.170 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2481.940 2658.170 2483.540 2738.170 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2328.340 2658.170 2329.940 2738.170 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2174.740 2658.170 2176.340 2738.170 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.140 2658.170 2022.740 2738.170 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2635.540 2145.030 2637.140 2225.030 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2481.940 2145.030 2483.540 2225.030 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2328.340 2145.030 2329.940 2225.030 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2174.740 2145.030 2176.340 2225.030 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.140 2145.030 2022.740 2225.030 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2635.540 1631.890 2637.140 1711.890 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2481.940 1631.890 2483.540 1711.890 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2328.340 1631.890 2329.940 1711.890 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2174.740 1631.890 2176.340 1711.890 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.140 1631.890 2022.740 1711.890 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2635.540 1118.750 2637.140 1198.750 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2481.940 1118.750 2483.540 1198.750 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2328.340 1118.750 2329.940 1198.750 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2174.740 1118.750 2176.340 1198.750 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.140 1118.750 2022.740 1198.750 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2635.540 605.610 2637.140 685.610 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2481.940 605.610 2483.540 685.610 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2328.340 605.610 2329.940 685.610 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2174.740 605.610 2176.340 685.610 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.140 605.610 2022.740 685.610 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2635.540 10.880 2637.140 172.470 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2481.940 10.880 2483.540 172.470 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2328.340 10.880 2329.940 172.470 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2174.740 10.880 2176.340 172.470 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.140 10.880 2022.740 172.470 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2558.740 3171.310 2560.340 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2405.140 3171.310 2406.740 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2251.540 3171.310 2253.140 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.940 3171.310 2099.540 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1944.340 10.880 1945.940 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1790.740 10.880 1792.340 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1637.140 10.880 1638.740 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1483.540 10.880 1485.140 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1329.940 10.880 1331.540 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1176.340 10.880 1177.940 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1022.740 10.880 1024.340 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.140 10.880 870.740 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2558.740 2658.170 2560.340 2738.170 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2405.140 2658.170 2406.740 2738.170 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2251.540 2658.170 2253.140 2738.170 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.940 2658.170 2099.540 2738.170 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2558.740 2145.030 2560.340 2225.030 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2405.140 2145.030 2406.740 2225.030 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2251.540 2145.030 2253.140 2225.030 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.940 2145.030 2099.540 2225.030 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2558.740 1631.890 2560.340 1711.890 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2405.140 1631.890 2406.740 1711.890 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2251.540 1631.890 2253.140 1711.890 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.940 1631.890 2099.540 1711.890 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2558.740 1118.750 2560.340 1198.750 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2405.140 1118.750 2406.740 1198.750 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2251.540 1118.750 2253.140 1198.750 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.940 1118.750 2099.540 1198.750 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2558.740 605.610 2560.340 685.610 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2405.140 605.610 2406.740 685.610 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2251.540 605.610 2253.140 685.610 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.940 605.610 2099.540 685.610 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2558.740 10.880 2560.340 172.470 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2405.140 10.880 2406.740 172.470 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2251.540 10.880 2253.140 172.470 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.940 10.880 2099.540 172.470 ;
    END
  END vssd2
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 2694.220 3288.565 ;
      LAYER met1 ;
        RECT 5.520 6.840 2699.670 3288.720 ;
      LAYER met2 ;
        RECT 5.680 3295.720 95.950 3296.000 ;
        RECT 96.790 3295.720 288.690 3296.000 ;
        RECT 289.530 3295.720 481.430 3296.000 ;
        RECT 482.270 3295.720 674.170 3296.000 ;
        RECT 675.010 3295.720 867.370 3296.000 ;
        RECT 868.210 3295.720 1060.110 3296.000 ;
        RECT 1060.950 3295.720 1252.850 3296.000 ;
        RECT 1253.690 3295.720 1446.050 3296.000 ;
        RECT 1446.890 3295.720 1638.790 3296.000 ;
        RECT 1639.630 3295.720 1831.530 3296.000 ;
        RECT 1832.370 3295.720 2024.270 3296.000 ;
        RECT 2025.110 3295.720 2217.470 3296.000 ;
        RECT 2218.310 3295.720 2410.210 3296.000 ;
        RECT 2411.050 3295.720 2602.950 3296.000 ;
        RECT 2603.790 3295.720 2699.640 3296.000 ;
        RECT 5.680 4.280 2699.640 3295.720 ;
        RECT 6.170 4.000 16.370 4.280 ;
        RECT 17.210 4.000 27.410 4.280 ;
        RECT 28.250 4.000 38.450 4.280 ;
        RECT 39.290 4.000 49.950 4.280 ;
        RECT 50.790 4.000 60.990 4.280 ;
        RECT 61.830 4.000 72.030 4.280 ;
        RECT 72.870 4.000 83.070 4.280 ;
        RECT 83.910 4.000 94.570 4.280 ;
        RECT 95.410 4.000 105.610 4.280 ;
        RECT 106.450 4.000 116.650 4.280 ;
        RECT 117.490 4.000 127.690 4.280 ;
        RECT 128.530 4.000 139.190 4.280 ;
        RECT 140.030 4.000 150.230 4.280 ;
        RECT 151.070 4.000 161.270 4.280 ;
        RECT 162.110 4.000 172.310 4.280 ;
        RECT 173.150 4.000 183.810 4.280 ;
        RECT 184.650 4.000 194.850 4.280 ;
        RECT 195.690 4.000 205.890 4.280 ;
        RECT 206.730 4.000 216.930 4.280 ;
        RECT 217.770 4.000 228.430 4.280 ;
        RECT 229.270 4.000 239.470 4.280 ;
        RECT 240.310 4.000 250.510 4.280 ;
        RECT 251.350 4.000 261.550 4.280 ;
        RECT 262.390 4.000 273.050 4.280 ;
        RECT 273.890 4.000 284.090 4.280 ;
        RECT 284.930 4.000 295.130 4.280 ;
        RECT 295.970 4.000 306.170 4.280 ;
        RECT 307.010 4.000 317.670 4.280 ;
        RECT 318.510 4.000 328.710 4.280 ;
        RECT 329.550 4.000 339.750 4.280 ;
        RECT 340.590 4.000 350.790 4.280 ;
        RECT 351.630 4.000 362.290 4.280 ;
        RECT 363.130 4.000 373.330 4.280 ;
        RECT 374.170 4.000 384.370 4.280 ;
        RECT 385.210 4.000 395.410 4.280 ;
        RECT 396.250 4.000 406.910 4.280 ;
        RECT 407.750 4.000 417.950 4.280 ;
        RECT 418.790 4.000 428.990 4.280 ;
        RECT 429.830 4.000 440.030 4.280 ;
        RECT 440.870 4.000 451.530 4.280 ;
        RECT 452.370 4.000 462.570 4.280 ;
        RECT 463.410 4.000 473.610 4.280 ;
        RECT 474.450 4.000 485.110 4.280 ;
        RECT 485.950 4.000 496.150 4.280 ;
        RECT 496.990 4.000 507.190 4.280 ;
        RECT 508.030 4.000 518.230 4.280 ;
        RECT 519.070 4.000 529.730 4.280 ;
        RECT 530.570 4.000 540.770 4.280 ;
        RECT 541.610 4.000 551.810 4.280 ;
        RECT 552.650 4.000 562.850 4.280 ;
        RECT 563.690 4.000 574.350 4.280 ;
        RECT 575.190 4.000 585.390 4.280 ;
        RECT 586.230 4.000 596.430 4.280 ;
        RECT 597.270 4.000 607.470 4.280 ;
        RECT 608.310 4.000 618.970 4.280 ;
        RECT 619.810 4.000 630.010 4.280 ;
        RECT 630.850 4.000 641.050 4.280 ;
        RECT 641.890 4.000 652.090 4.280 ;
        RECT 652.930 4.000 663.590 4.280 ;
        RECT 664.430 4.000 674.630 4.280 ;
        RECT 675.470 4.000 685.670 4.280 ;
        RECT 686.510 4.000 696.710 4.280 ;
        RECT 697.550 4.000 708.210 4.280 ;
        RECT 709.050 4.000 719.250 4.280 ;
        RECT 720.090 4.000 730.290 4.280 ;
        RECT 731.130 4.000 741.330 4.280 ;
        RECT 742.170 4.000 752.830 4.280 ;
        RECT 753.670 4.000 763.870 4.280 ;
        RECT 764.710 4.000 774.910 4.280 ;
        RECT 775.750 4.000 785.950 4.280 ;
        RECT 786.790 4.000 797.450 4.280 ;
        RECT 798.290 4.000 808.490 4.280 ;
        RECT 809.330 4.000 819.530 4.280 ;
        RECT 820.370 4.000 830.570 4.280 ;
        RECT 831.410 4.000 842.070 4.280 ;
        RECT 842.910 4.000 853.110 4.280 ;
        RECT 853.950 4.000 864.150 4.280 ;
        RECT 864.990 4.000 875.190 4.280 ;
        RECT 876.030 4.000 886.690 4.280 ;
        RECT 887.530 4.000 897.730 4.280 ;
        RECT 898.570 4.000 908.770 4.280 ;
        RECT 909.610 4.000 920.270 4.280 ;
        RECT 921.110 4.000 931.310 4.280 ;
        RECT 932.150 4.000 942.350 4.280 ;
        RECT 943.190 4.000 953.390 4.280 ;
        RECT 954.230 4.000 964.890 4.280 ;
        RECT 965.730 4.000 975.930 4.280 ;
        RECT 976.770 4.000 986.970 4.280 ;
        RECT 987.810 4.000 998.010 4.280 ;
        RECT 998.850 4.000 1009.510 4.280 ;
        RECT 1010.350 4.000 1020.550 4.280 ;
        RECT 1021.390 4.000 1031.590 4.280 ;
        RECT 1032.430 4.000 1042.630 4.280 ;
        RECT 1043.470 4.000 1054.130 4.280 ;
        RECT 1054.970 4.000 1065.170 4.280 ;
        RECT 1066.010 4.000 1076.210 4.280 ;
        RECT 1077.050 4.000 1087.250 4.280 ;
        RECT 1088.090 4.000 1098.750 4.280 ;
        RECT 1099.590 4.000 1109.790 4.280 ;
        RECT 1110.630 4.000 1120.830 4.280 ;
        RECT 1121.670 4.000 1131.870 4.280 ;
        RECT 1132.710 4.000 1143.370 4.280 ;
        RECT 1144.210 4.000 1154.410 4.280 ;
        RECT 1155.250 4.000 1165.450 4.280 ;
        RECT 1166.290 4.000 1176.490 4.280 ;
        RECT 1177.330 4.000 1187.990 4.280 ;
        RECT 1188.830 4.000 1199.030 4.280 ;
        RECT 1199.870 4.000 1210.070 4.280 ;
        RECT 1210.910 4.000 1221.110 4.280 ;
        RECT 1221.950 4.000 1232.610 4.280 ;
        RECT 1233.450 4.000 1243.650 4.280 ;
        RECT 1244.490 4.000 1254.690 4.280 ;
        RECT 1255.530 4.000 1265.730 4.280 ;
        RECT 1266.570 4.000 1277.230 4.280 ;
        RECT 1278.070 4.000 1288.270 4.280 ;
        RECT 1289.110 4.000 1299.310 4.280 ;
        RECT 1300.150 4.000 1310.350 4.280 ;
        RECT 1311.190 4.000 1321.850 4.280 ;
        RECT 1322.690 4.000 1332.890 4.280 ;
        RECT 1333.730 4.000 1343.930 4.280 ;
        RECT 1344.770 4.000 1355.430 4.280 ;
        RECT 1356.270 4.000 1366.470 4.280 ;
        RECT 1367.310 4.000 1377.510 4.280 ;
        RECT 1378.350 4.000 1388.550 4.280 ;
        RECT 1389.390 4.000 1400.050 4.280 ;
        RECT 1400.890 4.000 1411.090 4.280 ;
        RECT 1411.930 4.000 1422.130 4.280 ;
        RECT 1422.970 4.000 1433.170 4.280 ;
        RECT 1434.010 4.000 1444.670 4.280 ;
        RECT 1445.510 4.000 1455.710 4.280 ;
        RECT 1456.550 4.000 1466.750 4.280 ;
        RECT 1467.590 4.000 1477.790 4.280 ;
        RECT 1478.630 4.000 1489.290 4.280 ;
        RECT 1490.130 4.000 1500.330 4.280 ;
        RECT 1501.170 4.000 1511.370 4.280 ;
        RECT 1512.210 4.000 1522.410 4.280 ;
        RECT 1523.250 4.000 1533.910 4.280 ;
        RECT 1534.750 4.000 1544.950 4.280 ;
        RECT 1545.790 4.000 1555.990 4.280 ;
        RECT 1556.830 4.000 1567.030 4.280 ;
        RECT 1567.870 4.000 1578.530 4.280 ;
        RECT 1579.370 4.000 1589.570 4.280 ;
        RECT 1590.410 4.000 1600.610 4.280 ;
        RECT 1601.450 4.000 1611.650 4.280 ;
        RECT 1612.490 4.000 1623.150 4.280 ;
        RECT 1623.990 4.000 1634.190 4.280 ;
        RECT 1635.030 4.000 1645.230 4.280 ;
        RECT 1646.070 4.000 1656.270 4.280 ;
        RECT 1657.110 4.000 1667.770 4.280 ;
        RECT 1668.610 4.000 1678.810 4.280 ;
        RECT 1679.650 4.000 1689.850 4.280 ;
        RECT 1690.690 4.000 1700.890 4.280 ;
        RECT 1701.730 4.000 1712.390 4.280 ;
        RECT 1713.230 4.000 1723.430 4.280 ;
        RECT 1724.270 4.000 1734.470 4.280 ;
        RECT 1735.310 4.000 1745.510 4.280 ;
        RECT 1746.350 4.000 1757.010 4.280 ;
        RECT 1757.850 4.000 1768.050 4.280 ;
        RECT 1768.890 4.000 1779.090 4.280 ;
        RECT 1779.930 4.000 1790.130 4.280 ;
        RECT 1790.970 4.000 1801.630 4.280 ;
        RECT 1802.470 4.000 1812.670 4.280 ;
        RECT 1813.510 4.000 1823.710 4.280 ;
        RECT 1824.550 4.000 1835.210 4.280 ;
        RECT 1836.050 4.000 1846.250 4.280 ;
        RECT 1847.090 4.000 1857.290 4.280 ;
        RECT 1858.130 4.000 1868.330 4.280 ;
        RECT 1869.170 4.000 1879.830 4.280 ;
        RECT 1880.670 4.000 1890.870 4.280 ;
        RECT 1891.710 4.000 1901.910 4.280 ;
        RECT 1902.750 4.000 1912.950 4.280 ;
        RECT 1913.790 4.000 1924.450 4.280 ;
        RECT 1925.290 4.000 1935.490 4.280 ;
        RECT 1936.330 4.000 1946.530 4.280 ;
        RECT 1947.370 4.000 1957.570 4.280 ;
        RECT 1958.410 4.000 1969.070 4.280 ;
        RECT 1969.910 4.000 1980.110 4.280 ;
        RECT 1980.950 4.000 1991.150 4.280 ;
        RECT 1991.990 4.000 2002.190 4.280 ;
        RECT 2003.030 4.000 2013.690 4.280 ;
        RECT 2014.530 4.000 2024.730 4.280 ;
        RECT 2025.570 4.000 2035.770 4.280 ;
        RECT 2036.610 4.000 2046.810 4.280 ;
        RECT 2047.650 4.000 2058.310 4.280 ;
        RECT 2059.150 4.000 2069.350 4.280 ;
        RECT 2070.190 4.000 2080.390 4.280 ;
        RECT 2081.230 4.000 2091.430 4.280 ;
        RECT 2092.270 4.000 2102.930 4.280 ;
        RECT 2103.770 4.000 2113.970 4.280 ;
        RECT 2114.810 4.000 2125.010 4.280 ;
        RECT 2125.850 4.000 2136.050 4.280 ;
        RECT 2136.890 4.000 2147.550 4.280 ;
        RECT 2148.390 4.000 2158.590 4.280 ;
        RECT 2159.430 4.000 2169.630 4.280 ;
        RECT 2170.470 4.000 2180.670 4.280 ;
        RECT 2181.510 4.000 2192.170 4.280 ;
        RECT 2193.010 4.000 2203.210 4.280 ;
        RECT 2204.050 4.000 2214.250 4.280 ;
        RECT 2215.090 4.000 2225.290 4.280 ;
        RECT 2226.130 4.000 2236.790 4.280 ;
        RECT 2237.630 4.000 2247.830 4.280 ;
        RECT 2248.670 4.000 2258.870 4.280 ;
        RECT 2259.710 4.000 2270.370 4.280 ;
        RECT 2271.210 4.000 2281.410 4.280 ;
        RECT 2282.250 4.000 2292.450 4.280 ;
        RECT 2293.290 4.000 2303.490 4.280 ;
        RECT 2304.330 4.000 2314.990 4.280 ;
        RECT 2315.830 4.000 2326.030 4.280 ;
        RECT 2326.870 4.000 2337.070 4.280 ;
        RECT 2337.910 4.000 2348.110 4.280 ;
        RECT 2348.950 4.000 2359.610 4.280 ;
        RECT 2360.450 4.000 2370.650 4.280 ;
        RECT 2371.490 4.000 2381.690 4.280 ;
        RECT 2382.530 4.000 2392.730 4.280 ;
        RECT 2393.570 4.000 2404.230 4.280 ;
        RECT 2405.070 4.000 2415.270 4.280 ;
        RECT 2416.110 4.000 2426.310 4.280 ;
        RECT 2427.150 4.000 2437.350 4.280 ;
        RECT 2438.190 4.000 2448.850 4.280 ;
        RECT 2449.690 4.000 2459.890 4.280 ;
        RECT 2460.730 4.000 2470.930 4.280 ;
        RECT 2471.770 4.000 2481.970 4.280 ;
        RECT 2482.810 4.000 2493.470 4.280 ;
        RECT 2494.310 4.000 2504.510 4.280 ;
        RECT 2505.350 4.000 2515.550 4.280 ;
        RECT 2516.390 4.000 2526.590 4.280 ;
        RECT 2527.430 4.000 2538.090 4.280 ;
        RECT 2538.930 4.000 2549.130 4.280 ;
        RECT 2549.970 4.000 2560.170 4.280 ;
        RECT 2561.010 4.000 2571.210 4.280 ;
        RECT 2572.050 4.000 2582.710 4.280 ;
        RECT 2583.550 4.000 2593.750 4.280 ;
        RECT 2594.590 4.000 2604.790 4.280 ;
        RECT 2605.630 4.000 2615.830 4.280 ;
        RECT 2616.670 4.000 2627.330 4.280 ;
        RECT 2628.170 4.000 2638.370 4.280 ;
        RECT 2639.210 4.000 2649.410 4.280 ;
        RECT 2650.250 4.000 2660.450 4.280 ;
        RECT 2661.290 4.000 2671.950 4.280 ;
        RECT 2672.790 4.000 2682.990 4.280 ;
        RECT 2683.830 4.000 2694.030 4.280 ;
        RECT 2694.870 4.000 2699.640 4.280 ;
      LAYER met3 ;
        RECT 4.000 3150.120 2696.455 3288.645 ;
        RECT 4.400 3148.720 2696.455 3150.120 ;
        RECT 4.000 3025.680 2696.455 3148.720 ;
        RECT 4.000 3024.280 2695.600 3025.680 ;
        RECT 4.000 2850.240 2696.455 3024.280 ;
        RECT 4.400 2848.840 2696.455 2850.240 ;
        RECT 4.000 2550.360 2696.455 2848.840 ;
        RECT 4.400 2548.960 2696.455 2550.360 ;
        RECT 4.000 2475.560 2696.455 2548.960 ;
        RECT 4.000 2474.160 2695.600 2475.560 ;
        RECT 4.000 2250.480 2696.455 2474.160 ;
        RECT 4.400 2249.080 2696.455 2250.480 ;
        RECT 4.000 1950.600 2696.455 2249.080 ;
        RECT 4.400 1949.200 2696.455 1950.600 ;
        RECT 4.000 1925.440 2696.455 1949.200 ;
        RECT 4.000 1924.040 2695.600 1925.440 ;
        RECT 4.000 1650.040 2696.455 1924.040 ;
        RECT 4.400 1648.640 2696.455 1650.040 ;
        RECT 4.000 1375.320 2696.455 1648.640 ;
        RECT 4.000 1373.920 2695.600 1375.320 ;
        RECT 4.000 1350.160 2696.455 1373.920 ;
        RECT 4.400 1348.760 2696.455 1350.160 ;
        RECT 4.000 1050.280 2696.455 1348.760 ;
        RECT 4.400 1048.880 2696.455 1050.280 ;
        RECT 4.000 825.200 2696.455 1048.880 ;
        RECT 4.000 823.800 2695.600 825.200 ;
        RECT 4.000 750.400 2696.455 823.800 ;
        RECT 4.400 749.000 2696.455 750.400 ;
        RECT 4.000 450.520 2696.455 749.000 ;
        RECT 4.400 449.120 2696.455 450.520 ;
        RECT 4.000 275.760 2696.455 449.120 ;
        RECT 4.000 274.360 2695.600 275.760 ;
        RECT 4.000 150.640 2696.455 274.360 ;
        RECT 4.400 149.240 2696.455 150.640 ;
        RECT 4.000 10.715 2696.455 149.240 ;
      LAYER met4 ;
        RECT 432.695 17.175 481.440 3174.745 ;
        RECT 483.840 17.175 484.740 3174.745 ;
        RECT 487.140 17.175 558.240 3174.745 ;
        RECT 560.640 17.175 561.540 3174.745 ;
        RECT 563.940 17.175 635.040 3174.745 ;
        RECT 637.440 17.175 638.340 3174.745 ;
        RECT 640.740 17.175 711.840 3174.745 ;
        RECT 714.240 17.175 715.140 3174.745 ;
        RECT 717.540 17.175 788.640 3174.745 ;
        RECT 791.040 17.175 791.940 3174.745 ;
        RECT 794.340 17.175 865.440 3174.745 ;
        RECT 867.840 17.175 868.740 3174.745 ;
        RECT 871.140 17.175 942.240 3174.745 ;
        RECT 944.640 17.175 945.540 3174.745 ;
        RECT 947.940 17.175 1019.040 3174.745 ;
        RECT 1021.440 17.175 1022.340 3174.745 ;
        RECT 1024.740 17.175 1095.840 3174.745 ;
        RECT 1098.240 17.175 1099.140 3174.745 ;
        RECT 1101.540 17.175 1172.640 3174.745 ;
        RECT 1175.040 17.175 1175.940 3174.745 ;
        RECT 1178.340 17.175 1249.440 3174.745 ;
        RECT 1251.840 17.175 1252.740 3174.745 ;
        RECT 1255.140 17.175 1326.240 3174.745 ;
        RECT 1328.640 17.175 1329.540 3174.745 ;
        RECT 1331.940 17.175 1403.040 3174.745 ;
        RECT 1405.440 17.175 1406.340 3174.745 ;
        RECT 1408.740 17.175 1479.840 3174.745 ;
        RECT 1482.240 17.175 1483.140 3174.745 ;
        RECT 1485.540 17.175 1556.640 3174.745 ;
        RECT 1559.040 17.175 1559.940 3174.745 ;
        RECT 1562.340 17.175 1633.440 3174.745 ;
        RECT 1635.840 17.175 1636.740 3174.745 ;
        RECT 1639.140 17.175 1710.240 3174.745 ;
        RECT 1712.640 17.175 1713.540 3174.745 ;
        RECT 1715.940 17.175 1787.040 3174.745 ;
        RECT 1789.440 17.175 1790.340 3174.745 ;
        RECT 1792.740 17.175 1863.840 3174.745 ;
        RECT 1866.240 17.175 1867.140 3174.745 ;
        RECT 1869.540 17.175 1940.640 3174.745 ;
        RECT 1943.040 17.175 1943.940 3174.745 ;
        RECT 1946.340 3170.670 2017.440 3174.745 ;
        RECT 2019.840 3170.910 2020.740 3174.745 ;
        RECT 2023.140 3170.910 2094.240 3174.745 ;
        RECT 2019.840 3170.670 2094.240 3170.910 ;
        RECT 2096.640 3170.910 2097.540 3174.745 ;
        RECT 2099.940 3170.910 2171.040 3174.745 ;
        RECT 2096.640 3170.670 2171.040 3170.910 ;
        RECT 2173.440 3170.910 2174.340 3174.745 ;
        RECT 2176.740 3170.910 2247.840 3174.745 ;
        RECT 2173.440 3170.670 2247.840 3170.910 ;
        RECT 2250.240 3170.910 2251.140 3174.745 ;
        RECT 2253.540 3170.910 2324.640 3174.745 ;
        RECT 2250.240 3170.670 2324.640 3170.910 ;
        RECT 2327.040 3170.910 2327.940 3174.745 ;
        RECT 2330.340 3170.910 2401.440 3174.745 ;
        RECT 2327.040 3170.670 2401.440 3170.910 ;
        RECT 2403.840 3170.910 2404.740 3174.745 ;
        RECT 2407.140 3170.910 2478.240 3174.745 ;
        RECT 2403.840 3170.670 2478.240 3170.910 ;
        RECT 2480.640 3170.910 2481.540 3174.745 ;
        RECT 2483.940 3170.910 2555.040 3174.745 ;
        RECT 2480.640 3170.670 2555.040 3170.910 ;
        RECT 2557.440 3170.910 2558.340 3174.745 ;
        RECT 2560.740 3170.910 2631.840 3174.745 ;
        RECT 2557.440 3170.670 2631.840 3170.910 ;
        RECT 2634.240 3170.910 2635.140 3174.745 ;
        RECT 2637.540 3170.910 2693.465 3174.745 ;
        RECT 2634.240 3170.670 2693.465 3170.910 ;
        RECT 1946.340 2738.810 2693.465 3170.670 ;
        RECT 1946.340 2657.530 2017.440 2738.810 ;
        RECT 2019.840 2738.570 2094.240 2738.810 ;
        RECT 2019.840 2657.770 2020.740 2738.570 ;
        RECT 2023.140 2657.770 2094.240 2738.570 ;
        RECT 2019.840 2657.530 2094.240 2657.770 ;
        RECT 2096.640 2738.570 2171.040 2738.810 ;
        RECT 2096.640 2657.770 2097.540 2738.570 ;
        RECT 2099.940 2657.770 2171.040 2738.570 ;
        RECT 2096.640 2657.530 2171.040 2657.770 ;
        RECT 2173.440 2738.570 2247.840 2738.810 ;
        RECT 2173.440 2657.770 2174.340 2738.570 ;
        RECT 2176.740 2657.770 2247.840 2738.570 ;
        RECT 2173.440 2657.530 2247.840 2657.770 ;
        RECT 2250.240 2738.570 2324.640 2738.810 ;
        RECT 2250.240 2657.770 2251.140 2738.570 ;
        RECT 2253.540 2657.770 2324.640 2738.570 ;
        RECT 2250.240 2657.530 2324.640 2657.770 ;
        RECT 2327.040 2738.570 2401.440 2738.810 ;
        RECT 2327.040 2657.770 2327.940 2738.570 ;
        RECT 2330.340 2657.770 2401.440 2738.570 ;
        RECT 2327.040 2657.530 2401.440 2657.770 ;
        RECT 2403.840 2738.570 2478.240 2738.810 ;
        RECT 2403.840 2657.770 2404.740 2738.570 ;
        RECT 2407.140 2657.770 2478.240 2738.570 ;
        RECT 2403.840 2657.530 2478.240 2657.770 ;
        RECT 2480.640 2738.570 2555.040 2738.810 ;
        RECT 2480.640 2657.770 2481.540 2738.570 ;
        RECT 2483.940 2657.770 2555.040 2738.570 ;
        RECT 2480.640 2657.530 2555.040 2657.770 ;
        RECT 2557.440 2738.570 2631.840 2738.810 ;
        RECT 2557.440 2657.770 2558.340 2738.570 ;
        RECT 2560.740 2657.770 2631.840 2738.570 ;
        RECT 2557.440 2657.530 2631.840 2657.770 ;
        RECT 2634.240 2738.570 2693.465 2738.810 ;
        RECT 2634.240 2657.770 2635.140 2738.570 ;
        RECT 2637.540 2657.770 2693.465 2738.570 ;
        RECT 2634.240 2657.530 2693.465 2657.770 ;
        RECT 1946.340 2225.670 2693.465 2657.530 ;
        RECT 1946.340 2144.390 2017.440 2225.670 ;
        RECT 2019.840 2225.430 2094.240 2225.670 ;
        RECT 2019.840 2144.630 2020.740 2225.430 ;
        RECT 2023.140 2144.630 2094.240 2225.430 ;
        RECT 2019.840 2144.390 2094.240 2144.630 ;
        RECT 2096.640 2225.430 2171.040 2225.670 ;
        RECT 2096.640 2144.630 2097.540 2225.430 ;
        RECT 2099.940 2144.630 2171.040 2225.430 ;
        RECT 2096.640 2144.390 2171.040 2144.630 ;
        RECT 2173.440 2225.430 2247.840 2225.670 ;
        RECT 2173.440 2144.630 2174.340 2225.430 ;
        RECT 2176.740 2144.630 2247.840 2225.430 ;
        RECT 2173.440 2144.390 2247.840 2144.630 ;
        RECT 2250.240 2225.430 2324.640 2225.670 ;
        RECT 2250.240 2144.630 2251.140 2225.430 ;
        RECT 2253.540 2144.630 2324.640 2225.430 ;
        RECT 2250.240 2144.390 2324.640 2144.630 ;
        RECT 2327.040 2225.430 2401.440 2225.670 ;
        RECT 2327.040 2144.630 2327.940 2225.430 ;
        RECT 2330.340 2144.630 2401.440 2225.430 ;
        RECT 2327.040 2144.390 2401.440 2144.630 ;
        RECT 2403.840 2225.430 2478.240 2225.670 ;
        RECT 2403.840 2144.630 2404.740 2225.430 ;
        RECT 2407.140 2144.630 2478.240 2225.430 ;
        RECT 2403.840 2144.390 2478.240 2144.630 ;
        RECT 2480.640 2225.430 2555.040 2225.670 ;
        RECT 2480.640 2144.630 2481.540 2225.430 ;
        RECT 2483.940 2144.630 2555.040 2225.430 ;
        RECT 2480.640 2144.390 2555.040 2144.630 ;
        RECT 2557.440 2225.430 2631.840 2225.670 ;
        RECT 2557.440 2144.630 2558.340 2225.430 ;
        RECT 2560.740 2144.630 2631.840 2225.430 ;
        RECT 2557.440 2144.390 2631.840 2144.630 ;
        RECT 2634.240 2225.430 2693.465 2225.670 ;
        RECT 2634.240 2144.630 2635.140 2225.430 ;
        RECT 2637.540 2144.630 2693.465 2225.430 ;
        RECT 2634.240 2144.390 2693.465 2144.630 ;
        RECT 1946.340 1712.530 2693.465 2144.390 ;
        RECT 1946.340 1631.250 2017.440 1712.530 ;
        RECT 2019.840 1712.290 2094.240 1712.530 ;
        RECT 2019.840 1631.490 2020.740 1712.290 ;
        RECT 2023.140 1631.490 2094.240 1712.290 ;
        RECT 2019.840 1631.250 2094.240 1631.490 ;
        RECT 2096.640 1712.290 2171.040 1712.530 ;
        RECT 2096.640 1631.490 2097.540 1712.290 ;
        RECT 2099.940 1631.490 2171.040 1712.290 ;
        RECT 2096.640 1631.250 2171.040 1631.490 ;
        RECT 2173.440 1712.290 2247.840 1712.530 ;
        RECT 2173.440 1631.490 2174.340 1712.290 ;
        RECT 2176.740 1631.490 2247.840 1712.290 ;
        RECT 2173.440 1631.250 2247.840 1631.490 ;
        RECT 2250.240 1712.290 2324.640 1712.530 ;
        RECT 2250.240 1631.490 2251.140 1712.290 ;
        RECT 2253.540 1631.490 2324.640 1712.290 ;
        RECT 2250.240 1631.250 2324.640 1631.490 ;
        RECT 2327.040 1712.290 2401.440 1712.530 ;
        RECT 2327.040 1631.490 2327.940 1712.290 ;
        RECT 2330.340 1631.490 2401.440 1712.290 ;
        RECT 2327.040 1631.250 2401.440 1631.490 ;
        RECT 2403.840 1712.290 2478.240 1712.530 ;
        RECT 2403.840 1631.490 2404.740 1712.290 ;
        RECT 2407.140 1631.490 2478.240 1712.290 ;
        RECT 2403.840 1631.250 2478.240 1631.490 ;
        RECT 2480.640 1712.290 2555.040 1712.530 ;
        RECT 2480.640 1631.490 2481.540 1712.290 ;
        RECT 2483.940 1631.490 2555.040 1712.290 ;
        RECT 2480.640 1631.250 2555.040 1631.490 ;
        RECT 2557.440 1712.290 2631.840 1712.530 ;
        RECT 2557.440 1631.490 2558.340 1712.290 ;
        RECT 2560.740 1631.490 2631.840 1712.290 ;
        RECT 2557.440 1631.250 2631.840 1631.490 ;
        RECT 2634.240 1712.290 2693.465 1712.530 ;
        RECT 2634.240 1631.490 2635.140 1712.290 ;
        RECT 2637.540 1631.490 2693.465 1712.290 ;
        RECT 2634.240 1631.250 2693.465 1631.490 ;
        RECT 1946.340 1199.390 2693.465 1631.250 ;
        RECT 1946.340 1118.110 2017.440 1199.390 ;
        RECT 2019.840 1199.150 2094.240 1199.390 ;
        RECT 2019.840 1118.350 2020.740 1199.150 ;
        RECT 2023.140 1118.350 2094.240 1199.150 ;
        RECT 2019.840 1118.110 2094.240 1118.350 ;
        RECT 2096.640 1199.150 2171.040 1199.390 ;
        RECT 2096.640 1118.350 2097.540 1199.150 ;
        RECT 2099.940 1118.350 2171.040 1199.150 ;
        RECT 2096.640 1118.110 2171.040 1118.350 ;
        RECT 2173.440 1199.150 2247.840 1199.390 ;
        RECT 2173.440 1118.350 2174.340 1199.150 ;
        RECT 2176.740 1118.350 2247.840 1199.150 ;
        RECT 2173.440 1118.110 2247.840 1118.350 ;
        RECT 2250.240 1199.150 2324.640 1199.390 ;
        RECT 2250.240 1118.350 2251.140 1199.150 ;
        RECT 2253.540 1118.350 2324.640 1199.150 ;
        RECT 2250.240 1118.110 2324.640 1118.350 ;
        RECT 2327.040 1199.150 2401.440 1199.390 ;
        RECT 2327.040 1118.350 2327.940 1199.150 ;
        RECT 2330.340 1118.350 2401.440 1199.150 ;
        RECT 2327.040 1118.110 2401.440 1118.350 ;
        RECT 2403.840 1199.150 2478.240 1199.390 ;
        RECT 2403.840 1118.350 2404.740 1199.150 ;
        RECT 2407.140 1118.350 2478.240 1199.150 ;
        RECT 2403.840 1118.110 2478.240 1118.350 ;
        RECT 2480.640 1199.150 2555.040 1199.390 ;
        RECT 2480.640 1118.350 2481.540 1199.150 ;
        RECT 2483.940 1118.350 2555.040 1199.150 ;
        RECT 2480.640 1118.110 2555.040 1118.350 ;
        RECT 2557.440 1199.150 2631.840 1199.390 ;
        RECT 2557.440 1118.350 2558.340 1199.150 ;
        RECT 2560.740 1118.350 2631.840 1199.150 ;
        RECT 2557.440 1118.110 2631.840 1118.350 ;
        RECT 2634.240 1199.150 2693.465 1199.390 ;
        RECT 2634.240 1118.350 2635.140 1199.150 ;
        RECT 2637.540 1118.350 2693.465 1199.150 ;
        RECT 2634.240 1118.110 2693.465 1118.350 ;
        RECT 1946.340 686.250 2693.465 1118.110 ;
        RECT 1946.340 604.970 2017.440 686.250 ;
        RECT 2019.840 686.010 2094.240 686.250 ;
        RECT 2019.840 605.210 2020.740 686.010 ;
        RECT 2023.140 605.210 2094.240 686.010 ;
        RECT 2019.840 604.970 2094.240 605.210 ;
        RECT 2096.640 686.010 2171.040 686.250 ;
        RECT 2096.640 605.210 2097.540 686.010 ;
        RECT 2099.940 605.210 2171.040 686.010 ;
        RECT 2096.640 604.970 2171.040 605.210 ;
        RECT 2173.440 686.010 2247.840 686.250 ;
        RECT 2173.440 605.210 2174.340 686.010 ;
        RECT 2176.740 605.210 2247.840 686.010 ;
        RECT 2173.440 604.970 2247.840 605.210 ;
        RECT 2250.240 686.010 2324.640 686.250 ;
        RECT 2250.240 605.210 2251.140 686.010 ;
        RECT 2253.540 605.210 2324.640 686.010 ;
        RECT 2250.240 604.970 2324.640 605.210 ;
        RECT 2327.040 686.010 2401.440 686.250 ;
        RECT 2327.040 605.210 2327.940 686.010 ;
        RECT 2330.340 605.210 2401.440 686.010 ;
        RECT 2327.040 604.970 2401.440 605.210 ;
        RECT 2403.840 686.010 2478.240 686.250 ;
        RECT 2403.840 605.210 2404.740 686.010 ;
        RECT 2407.140 605.210 2478.240 686.010 ;
        RECT 2403.840 604.970 2478.240 605.210 ;
        RECT 2480.640 686.010 2555.040 686.250 ;
        RECT 2480.640 605.210 2481.540 686.010 ;
        RECT 2483.940 605.210 2555.040 686.010 ;
        RECT 2480.640 604.970 2555.040 605.210 ;
        RECT 2557.440 686.010 2631.840 686.250 ;
        RECT 2557.440 605.210 2558.340 686.010 ;
        RECT 2560.740 605.210 2631.840 686.010 ;
        RECT 2557.440 604.970 2631.840 605.210 ;
        RECT 2634.240 686.010 2693.465 686.250 ;
        RECT 2634.240 605.210 2635.140 686.010 ;
        RECT 2637.540 605.210 2693.465 686.010 ;
        RECT 2634.240 604.970 2693.465 605.210 ;
        RECT 1946.340 173.110 2693.465 604.970 ;
        RECT 1946.340 17.175 2017.440 173.110 ;
        RECT 2019.840 172.870 2094.240 173.110 ;
        RECT 2019.840 17.175 2020.740 172.870 ;
        RECT 2023.140 17.175 2094.240 172.870 ;
        RECT 2096.640 172.870 2171.040 173.110 ;
        RECT 2096.640 17.175 2097.540 172.870 ;
        RECT 2099.940 17.175 2171.040 172.870 ;
        RECT 2173.440 172.870 2247.840 173.110 ;
        RECT 2173.440 17.175 2174.340 172.870 ;
        RECT 2176.740 17.175 2247.840 172.870 ;
        RECT 2250.240 172.870 2324.640 173.110 ;
        RECT 2250.240 17.175 2251.140 172.870 ;
        RECT 2253.540 17.175 2324.640 172.870 ;
        RECT 2327.040 172.870 2401.440 173.110 ;
        RECT 2327.040 17.175 2327.940 172.870 ;
        RECT 2330.340 17.175 2401.440 172.870 ;
        RECT 2403.840 172.870 2478.240 173.110 ;
        RECT 2403.840 17.175 2404.740 172.870 ;
        RECT 2407.140 17.175 2478.240 172.870 ;
        RECT 2480.640 172.870 2555.040 173.110 ;
        RECT 2480.640 17.175 2481.540 172.870 ;
        RECT 2483.940 17.175 2555.040 172.870 ;
        RECT 2557.440 172.870 2631.840 173.110 ;
        RECT 2557.440 17.175 2558.340 172.870 ;
        RECT 2560.740 17.175 2631.840 172.870 ;
        RECT 2634.240 172.870 2693.465 173.110 ;
        RECT 2634.240 17.175 2635.140 172.870 ;
        RECT 2637.540 17.175 2693.465 172.870 ;
  END
END top_level_bASIC
END LIBRARY


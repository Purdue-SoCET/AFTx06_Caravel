VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_level_bASIC
  CLASS BLOCK ;
  FOREIGN top_level_bASIC ;
  ORIGIN 0.000 0.000 ;
  SIZE 2700.000 BY 3300.000 ;
  PIN MISO_bi
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.190 3296.000 1350.470 3300.000 ;
    END
  END MISO_bi
  PIN MISO_output_en_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 3296.000 810.430 3300.000 ;
    END
  END MISO_output_en_low
  PIN MOSI_bi
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2430.270 3296.000 2430.550 3300.000 ;
    END
  END MOSI_bi
  PIN MOSI_output_en_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.230 3296.000 1890.510 3300.000 ;
    END
  END MOSI_output_en_low
  PIN SCK_bi
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3033.520 2700.000 3034.120 ;
    END
  END SCK_bi
  PIN SCK_output_en_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3139.600 2700.000 3140.200 ;
    END
  END SCK_output_en_low
  PIN SCL_bi
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2607.840 2700.000 2608.440 ;
    END
  END SCL_bi
  PIN SCL_output_en_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2713.920 2700.000 2714.520 ;
    END
  END SCL_output_en_low
  PIN SDA_bi
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2395.000 2700.000 2395.600 ;
    END
  END SDA_bi
  PIN SDA_output_en_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2501.080 2700.000 2501.680 ;
    END
  END SDA_output_en_low
  PIN SS_bi
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2820.680 2700.000 2821.280 ;
    END
  END SS_bi
  PIN SS_output_en_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2926.760 2700.000 2927.360 ;
    END
  END SS_output_en_low
  PIN asyncrst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 265.920 2700.000 266.520 ;
    END
  END asyncrst_n
  PIN clk_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 53.080 2700.000 53.680 ;
    END
  END clk_sel
  PIN gpio_bidir_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 372.000 2700.000 372.600 ;
    END
  END gpio_bidir_io[0]
  PIN gpio_bidir_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 584.840 2700.000 585.440 ;
    END
  END gpio_bidir_io[1]
  PIN gpio_bidir_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 797.680 2700.000 798.280 ;
    END
  END gpio_bidir_io[2]
  PIN gpio_bidir_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1010.520 2700.000 1011.120 ;
    END
  END gpio_bidir_io[3]
  PIN gpio_bidir_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1224.040 2700.000 1224.640 ;
    END
  END gpio_bidir_io[4]
  PIN gpio_bidir_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1436.880 2700.000 1437.480 ;
    END
  END gpio_bidir_io[5]
  PIN gpio_bidir_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1649.720 2700.000 1650.320 ;
    END
  END gpio_bidir_io[6]
  PIN gpio_bidir_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1862.560 2700.000 1863.160 ;
    END
  END gpio_bidir_io[7]
  PIN gpio_output_en_low[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 478.760 2700.000 479.360 ;
    END
  END gpio_output_en_low[0]
  PIN gpio_output_en_low[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 691.600 2700.000 692.200 ;
    END
  END gpio_output_en_low[1]
  PIN gpio_output_en_low[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 904.440 2700.000 905.040 ;
    END
  END gpio_output_en_low[2]
  PIN gpio_output_en_low[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1117.280 2700.000 1117.880 ;
    END
  END gpio_output_en_low[3]
  PIN gpio_output_en_low[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1330.120 2700.000 1330.720 ;
    END
  END gpio_output_en_low[4]
  PIN gpio_output_en_low[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1542.960 2700.000 1543.560 ;
    END
  END gpio_output_en_low[5]
  PIN gpio_output_en_low[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1755.800 2700.000 1756.400 ;
    END
  END gpio_output_en_low[6]
  PIN gpio_output_en_low[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 1968.640 2700.000 1969.240 ;
    END
  END gpio_output_en_low[7]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 3296.000 270.390 3300.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3246.360 2700.000 3246.960 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2694.310 0.000 2694.590 4.000 ;
    END
  END irq[2]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.170 0.000 1218.450 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2362.190 0.000 2362.470 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2373.690 0.000 2373.970 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2385.190 0.000 2385.470 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.690 0.000 2396.970 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.190 0.000 2408.470 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2419.690 0.000 2419.970 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.190 0.000 2431.470 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2442.230 0.000 2442.510 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2453.730 0.000 2454.010 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2465.230 0.000 2465.510 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.710 0.000 1332.990 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2476.730 0.000 2477.010 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2488.230 0.000 2488.510 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2499.730 0.000 2500.010 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2511.230 0.000 2511.510 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2522.730 0.000 2523.010 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2533.770 0.000 2534.050 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2545.270 0.000 2545.550 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.770 0.000 2557.050 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2568.270 0.000 2568.550 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.770 0.000 2580.050 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.210 0.000 1344.490 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.270 0.000 2591.550 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2602.770 0.000 2603.050 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2614.270 0.000 2614.550 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2625.310 0.000 2625.590 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2636.810 0.000 2637.090 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2648.310 0.000 2648.590 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2659.810 0.000 2660.090 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2671.310 0.000 2671.590 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 0.000 1355.990 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.750 0.000 1367.030 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.250 0.000 1378.530 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1389.750 0.000 1390.030 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.250 0.000 1401.530 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.750 0.000 1413.030 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1424.250 0.000 1424.530 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.750 0.000 1436.030 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.670 0.000 1229.950 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.790 0.000 1447.070 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.290 0.000 1458.570 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1469.790 0.000 1470.070 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 0.000 1481.570 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.790 0.000 1493.070 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1504.290 0.000 1504.570 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.790 0.000 1516.070 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.290 0.000 1527.570 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1538.330 0.000 1538.610 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1549.830 0.000 1550.110 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.170 0.000 1241.450 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.330 0.000 1561.610 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.830 0.000 1573.110 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 0.000 1584.610 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1595.830 0.000 1596.110 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.330 0.000 1607.610 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.830 0.000 1619.110 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.870 0.000 1630.150 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1641.370 0.000 1641.650 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1652.870 0.000 1653.150 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.370 0.000 1664.650 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 0.000 1252.950 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.870 0.000 1676.150 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.370 0.000 1687.650 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1698.870 0.000 1699.150 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.370 0.000 1710.650 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.410 0.000 1721.690 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.910 0.000 1733.190 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1744.410 0.000 1744.690 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1755.910 0.000 1756.190 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.410 0.000 1767.690 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1778.910 0.000 1779.190 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.170 0.000 1264.450 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.410 0.000 1790.690 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1801.910 0.000 1802.190 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.950 0.000 1813.230 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.450 0.000 1824.730 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.950 0.000 1836.230 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1847.450 0.000 1847.730 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.950 0.000 1859.230 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.450 0.000 1870.730 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.950 0.000 1882.230 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.450 0.000 1893.730 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.210 0.000 1275.490 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.490 0.000 1904.770 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.990 0.000 1916.270 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.490 0.000 1927.770 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.990 0.000 1939.270 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1950.490 0.000 1950.770 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.990 0.000 1962.270 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1973.490 0.000 1973.770 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1984.990 0.000 1985.270 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1996.030 0.000 1996.310 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2007.530 0.000 2007.810 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.710 0.000 1286.990 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.030 0.000 2019.310 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.530 0.000 2030.810 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.030 0.000 2042.310 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.530 0.000 2053.810 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.030 0.000 2065.310 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2076.070 0.000 2076.350 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2087.570 0.000 2087.850 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.070 0.000 2099.350 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2110.570 0.000 2110.850 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2122.070 0.000 2122.350 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.210 0.000 1298.490 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2133.570 0.000 2133.850 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2145.070 0.000 2145.350 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2156.570 0.000 2156.850 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2167.610 0.000 2167.890 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2179.110 0.000 2179.390 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2190.610 0.000 2190.890 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2202.110 0.000 2202.390 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.610 0.000 2213.890 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2225.110 0.000 2225.390 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.610 0.000 2236.890 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.710 0.000 1309.990 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.110 0.000 2248.390 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2259.150 0.000 2259.430 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2270.650 0.000 2270.930 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2282.150 0.000 2282.430 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2293.650 0.000 2293.930 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2305.150 0.000 2305.430 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2316.650 0.000 2316.930 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.150 0.000 2328.430 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2339.650 0.000 2339.930 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2350.690 0.000 2350.970 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1321.210 0.000 1321.490 4.000 ;
    END
  END la_data_out[9]
  PIN pwm_w_data_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2075.400 2700.000 2076.000 ;
    END
  END pwm_w_data_0
  PIN timer_bidir_0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2181.480 2700.000 2182.080 ;
    END
  END timer_bidir_0
  PIN timer_output_en_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 2288.240 2700.000 2288.840 ;
    END
  END timer_output_en_low
  PIN uart_debug_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1649.720 4.000 1650.320 ;
    END
  END uart_debug_rx
  PIN uart_debug_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 159.160 2700.000 159.760 ;
    END
  END uart_debug_tx
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2682.810 0.000 2683.090 4.000 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 0.000 600.670 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 0.000 635.170 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 0.000 669.210 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.430 0.000 703.710 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 0.000 737.750 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 0.000 772.250 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 0.000 806.750 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 0.000 875.290 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.050 0.000 909.330 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.050 0.000 978.330 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.090 0.000 1012.370 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 0.000 1046.870 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.090 0.000 1081.370 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.130 0.000 1115.410 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 0.000 1149.910 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.670 0.000 1183.950 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 0.000 543.630 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 0.000 577.670 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 0.000 749.250 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.470 0.000 783.750 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.510 0.000 817.790 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.010 0.000 852.290 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.510 0.000 886.790 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 0.000 920.830 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 0.000 955.330 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.550 0.000 989.830 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.590 0.000 1023.870 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.090 0.000 1058.370 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.130 0.000 1092.410 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.630 0.000 1126.910 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.130 0.000 1161.410 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.170 0.000 1195.450 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 0.000 554.670 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 0.000 623.670 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 0.000 657.710 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.930 0.000 692.210 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 0.000 726.250 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.470 0.000 760.750 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 0.000 795.250 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 0.000 829.290 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.510 0.000 863.790 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.010 0.000 898.290 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.050 0.000 932.330 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 0.000 966.830 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.590 0.000 1000.870 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.090 0.000 1035.370 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.590 0.000 1069.870 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.630 0.000 1103.910 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.130 0.000 1138.410 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.630 0.000 1172.910 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.670 0.000 1206.950 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 3159.510 2633.840 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 3159.510 2480.240 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 3159.510 2326.640 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 3159.510 2173.040 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 3159.510 2019.440 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 3288.720 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 2646.370 2633.840 2738.410 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 2646.370 2480.240 2738.410 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 2646.370 2326.640 2738.410 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 2646.370 2173.040 2738.410 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 2646.370 2019.440 2738.410 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 2133.230 2633.840 2225.270 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 2133.230 2480.240 2225.270 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 2133.230 2326.640 2225.270 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 2133.230 2173.040 2225.270 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 2133.230 2019.440 2225.270 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 1620.090 2633.840 1712.130 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 1620.090 2480.240 1712.130 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 1620.090 2326.640 1712.130 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 1620.090 2173.040 1712.130 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 1620.090 2019.440 1712.130 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 1106.950 2633.840 1198.990 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 1106.950 2480.240 1198.990 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 1106.950 2326.640 1198.990 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 1106.950 2173.040 1198.990 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 1106.950 2019.440 1198.990 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 593.810 2633.840 685.850 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 593.810 2480.240 685.850 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 593.810 2326.640 685.850 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 593.810 2173.040 685.850 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 593.810 2019.440 685.850 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 172.710 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 172.710 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 172.710 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 172.710 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 172.710 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 3159.510 2557.040 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 3159.510 2403.440 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 3159.510 2249.840 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 3159.510 2096.240 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 3288.720 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 2646.370 2557.040 2738.410 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 2646.370 2403.440 2738.410 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 2646.370 2249.840 2738.410 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 2646.370 2096.240 2738.410 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 2133.230 2557.040 2225.270 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 2133.230 2403.440 2225.270 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 2133.230 2249.840 2225.270 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 2133.230 2096.240 2225.270 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 1620.090 2557.040 1712.130 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 1620.090 2403.440 1712.130 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 1620.090 2249.840 1712.130 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 1620.090 2096.240 1712.130 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 1106.950 2557.040 1198.990 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 1106.950 2403.440 1198.990 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 1106.950 2249.840 1198.990 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 1106.950 2096.240 1198.990 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 593.810 2557.040 685.850 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 593.810 2403.440 685.850 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 593.810 2249.840 685.850 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 593.810 2096.240 685.850 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 172.710 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 172.710 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 172.710 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 172.710 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2635.540 3159.750 2637.140 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2481.940 3159.750 2483.540 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2328.340 3159.750 2329.940 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2174.740 3159.750 2176.340 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.140 3159.750 2022.740 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1867.540 10.880 1869.140 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1713.940 10.880 1715.540 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1560.340 10.880 1561.940 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1406.740 10.880 1408.340 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1253.140 10.880 1254.740 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1099.540 10.880 1101.140 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 945.940 10.880 947.540 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.340 10.880 793.940 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 3288.480 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2635.540 2646.610 2637.140 2738.170 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2481.940 2646.610 2483.540 2738.170 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2328.340 2646.610 2329.940 2738.170 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2174.740 2646.610 2176.340 2738.170 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.140 2646.610 2022.740 2738.170 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2635.540 2133.470 2637.140 2225.030 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2481.940 2133.470 2483.540 2225.030 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2328.340 2133.470 2329.940 2225.030 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2174.740 2133.470 2176.340 2225.030 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.140 2133.470 2022.740 2225.030 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2635.540 1620.330 2637.140 1711.890 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2481.940 1620.330 2483.540 1711.890 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2328.340 1620.330 2329.940 1711.890 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2174.740 1620.330 2176.340 1711.890 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.140 1620.330 2022.740 1711.890 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2635.540 1107.190 2637.140 1198.750 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2481.940 1107.190 2483.540 1198.750 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2328.340 1107.190 2329.940 1198.750 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2174.740 1107.190 2176.340 1198.750 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.140 1107.190 2022.740 1198.750 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2635.540 594.050 2637.140 685.610 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2481.940 594.050 2483.540 685.610 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2328.340 594.050 2329.940 685.610 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2174.740 594.050 2176.340 685.610 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.140 594.050 2022.740 685.610 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2635.540 10.880 2637.140 172.470 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2481.940 10.880 2483.540 172.470 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2328.340 10.880 2329.940 172.470 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2174.740 10.880 2176.340 172.470 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.140 10.880 2022.740 172.470 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2558.740 3159.750 2560.340 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2405.140 3159.750 2406.740 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2251.540 3159.750 2253.140 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.940 3159.750 2099.540 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1944.340 10.880 1945.940 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1790.740 10.880 1792.340 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1637.140 10.880 1638.740 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1483.540 10.880 1485.140 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1329.940 10.880 1331.540 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1176.340 10.880 1177.940 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1022.740 10.880 1024.340 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.140 10.880 870.740 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 3288.480 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2558.740 2646.610 2560.340 2738.170 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2405.140 2646.610 2406.740 2738.170 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2251.540 2646.610 2253.140 2738.170 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.940 2646.610 2099.540 2738.170 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2558.740 2133.470 2560.340 2225.030 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2405.140 2133.470 2406.740 2225.030 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2251.540 2133.470 2253.140 2225.030 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.940 2133.470 2099.540 2225.030 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2558.740 1620.330 2560.340 1711.890 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2405.140 1620.330 2406.740 1711.890 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2251.540 1620.330 2253.140 1711.890 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.940 1620.330 2099.540 1711.890 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2558.740 1107.190 2560.340 1198.750 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2405.140 1107.190 2406.740 1198.750 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2251.540 1107.190 2253.140 1198.750 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.940 1107.190 2099.540 1198.750 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2558.740 594.050 2560.340 685.610 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2405.140 594.050 2406.740 685.610 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2251.540 594.050 2253.140 685.610 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.940 594.050 2099.540 685.610 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2558.740 10.880 2560.340 172.470 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2405.140 10.880 2406.740 172.470 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2251.540 10.880 2253.140 172.470 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.940 10.880 2099.540 172.470 ;
    END
  END vssd2
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 2694.220 3288.565 ;
      LAYER met1 ;
        RECT 5.520 6.840 2697.830 3288.720 ;
      LAYER met2 ;
        RECT 5.620 3295.720 269.830 3296.000 ;
        RECT 270.670 3295.720 809.870 3296.000 ;
        RECT 810.710 3295.720 1349.910 3296.000 ;
        RECT 1350.750 3295.720 1889.950 3296.000 ;
        RECT 1890.790 3295.720 2429.990 3296.000 ;
        RECT 2430.830 3295.720 2697.800 3296.000 ;
        RECT 5.620 4.280 2697.800 3295.720 ;
        RECT 6.170 4.000 16.370 4.280 ;
        RECT 17.210 4.000 27.870 4.280 ;
        RECT 28.710 4.000 39.370 4.280 ;
        RECT 40.210 4.000 50.870 4.280 ;
        RECT 51.710 4.000 62.370 4.280 ;
        RECT 63.210 4.000 73.870 4.280 ;
        RECT 74.710 4.000 85.370 4.280 ;
        RECT 86.210 4.000 96.410 4.280 ;
        RECT 97.250 4.000 107.910 4.280 ;
        RECT 108.750 4.000 119.410 4.280 ;
        RECT 120.250 4.000 130.910 4.280 ;
        RECT 131.750 4.000 142.410 4.280 ;
        RECT 143.250 4.000 153.910 4.280 ;
        RECT 154.750 4.000 165.410 4.280 ;
        RECT 166.250 4.000 176.910 4.280 ;
        RECT 177.750 4.000 187.950 4.280 ;
        RECT 188.790 4.000 199.450 4.280 ;
        RECT 200.290 4.000 210.950 4.280 ;
        RECT 211.790 4.000 222.450 4.280 ;
        RECT 223.290 4.000 233.950 4.280 ;
        RECT 234.790 4.000 245.450 4.280 ;
        RECT 246.290 4.000 256.950 4.280 ;
        RECT 257.790 4.000 268.450 4.280 ;
        RECT 269.290 4.000 279.490 4.280 ;
        RECT 280.330 4.000 290.990 4.280 ;
        RECT 291.830 4.000 302.490 4.280 ;
        RECT 303.330 4.000 313.990 4.280 ;
        RECT 314.830 4.000 325.490 4.280 ;
        RECT 326.330 4.000 336.990 4.280 ;
        RECT 337.830 4.000 348.490 4.280 ;
        RECT 349.330 4.000 359.990 4.280 ;
        RECT 360.830 4.000 371.030 4.280 ;
        RECT 371.870 4.000 382.530 4.280 ;
        RECT 383.370 4.000 394.030 4.280 ;
        RECT 394.870 4.000 405.530 4.280 ;
        RECT 406.370 4.000 417.030 4.280 ;
        RECT 417.870 4.000 428.530 4.280 ;
        RECT 429.370 4.000 440.030 4.280 ;
        RECT 440.870 4.000 451.530 4.280 ;
        RECT 452.370 4.000 462.570 4.280 ;
        RECT 463.410 4.000 474.070 4.280 ;
        RECT 474.910 4.000 485.570 4.280 ;
        RECT 486.410 4.000 497.070 4.280 ;
        RECT 497.910 4.000 508.570 4.280 ;
        RECT 509.410 4.000 520.070 4.280 ;
        RECT 520.910 4.000 531.570 4.280 ;
        RECT 532.410 4.000 543.070 4.280 ;
        RECT 543.910 4.000 554.110 4.280 ;
        RECT 554.950 4.000 565.610 4.280 ;
        RECT 566.450 4.000 577.110 4.280 ;
        RECT 577.950 4.000 588.610 4.280 ;
        RECT 589.450 4.000 600.110 4.280 ;
        RECT 600.950 4.000 611.610 4.280 ;
        RECT 612.450 4.000 623.110 4.280 ;
        RECT 623.950 4.000 634.610 4.280 ;
        RECT 635.450 4.000 645.650 4.280 ;
        RECT 646.490 4.000 657.150 4.280 ;
        RECT 657.990 4.000 668.650 4.280 ;
        RECT 669.490 4.000 680.150 4.280 ;
        RECT 680.990 4.000 691.650 4.280 ;
        RECT 692.490 4.000 703.150 4.280 ;
        RECT 703.990 4.000 714.650 4.280 ;
        RECT 715.490 4.000 725.690 4.280 ;
        RECT 726.530 4.000 737.190 4.280 ;
        RECT 738.030 4.000 748.690 4.280 ;
        RECT 749.530 4.000 760.190 4.280 ;
        RECT 761.030 4.000 771.690 4.280 ;
        RECT 772.530 4.000 783.190 4.280 ;
        RECT 784.030 4.000 794.690 4.280 ;
        RECT 795.530 4.000 806.190 4.280 ;
        RECT 807.030 4.000 817.230 4.280 ;
        RECT 818.070 4.000 828.730 4.280 ;
        RECT 829.570 4.000 840.230 4.280 ;
        RECT 841.070 4.000 851.730 4.280 ;
        RECT 852.570 4.000 863.230 4.280 ;
        RECT 864.070 4.000 874.730 4.280 ;
        RECT 875.570 4.000 886.230 4.280 ;
        RECT 887.070 4.000 897.730 4.280 ;
        RECT 898.570 4.000 908.770 4.280 ;
        RECT 909.610 4.000 920.270 4.280 ;
        RECT 921.110 4.000 931.770 4.280 ;
        RECT 932.610 4.000 943.270 4.280 ;
        RECT 944.110 4.000 954.770 4.280 ;
        RECT 955.610 4.000 966.270 4.280 ;
        RECT 967.110 4.000 977.770 4.280 ;
        RECT 978.610 4.000 989.270 4.280 ;
        RECT 990.110 4.000 1000.310 4.280 ;
        RECT 1001.150 4.000 1011.810 4.280 ;
        RECT 1012.650 4.000 1023.310 4.280 ;
        RECT 1024.150 4.000 1034.810 4.280 ;
        RECT 1035.650 4.000 1046.310 4.280 ;
        RECT 1047.150 4.000 1057.810 4.280 ;
        RECT 1058.650 4.000 1069.310 4.280 ;
        RECT 1070.150 4.000 1080.810 4.280 ;
        RECT 1081.650 4.000 1091.850 4.280 ;
        RECT 1092.690 4.000 1103.350 4.280 ;
        RECT 1104.190 4.000 1114.850 4.280 ;
        RECT 1115.690 4.000 1126.350 4.280 ;
        RECT 1127.190 4.000 1137.850 4.280 ;
        RECT 1138.690 4.000 1149.350 4.280 ;
        RECT 1150.190 4.000 1160.850 4.280 ;
        RECT 1161.690 4.000 1172.350 4.280 ;
        RECT 1173.190 4.000 1183.390 4.280 ;
        RECT 1184.230 4.000 1194.890 4.280 ;
        RECT 1195.730 4.000 1206.390 4.280 ;
        RECT 1207.230 4.000 1217.890 4.280 ;
        RECT 1218.730 4.000 1229.390 4.280 ;
        RECT 1230.230 4.000 1240.890 4.280 ;
        RECT 1241.730 4.000 1252.390 4.280 ;
        RECT 1253.230 4.000 1263.890 4.280 ;
        RECT 1264.730 4.000 1274.930 4.280 ;
        RECT 1275.770 4.000 1286.430 4.280 ;
        RECT 1287.270 4.000 1297.930 4.280 ;
        RECT 1298.770 4.000 1309.430 4.280 ;
        RECT 1310.270 4.000 1320.930 4.280 ;
        RECT 1321.770 4.000 1332.430 4.280 ;
        RECT 1333.270 4.000 1343.930 4.280 ;
        RECT 1344.770 4.000 1355.430 4.280 ;
        RECT 1356.270 4.000 1366.470 4.280 ;
        RECT 1367.310 4.000 1377.970 4.280 ;
        RECT 1378.810 4.000 1389.470 4.280 ;
        RECT 1390.310 4.000 1400.970 4.280 ;
        RECT 1401.810 4.000 1412.470 4.280 ;
        RECT 1413.310 4.000 1423.970 4.280 ;
        RECT 1424.810 4.000 1435.470 4.280 ;
        RECT 1436.310 4.000 1446.510 4.280 ;
        RECT 1447.350 4.000 1458.010 4.280 ;
        RECT 1458.850 4.000 1469.510 4.280 ;
        RECT 1470.350 4.000 1481.010 4.280 ;
        RECT 1481.850 4.000 1492.510 4.280 ;
        RECT 1493.350 4.000 1504.010 4.280 ;
        RECT 1504.850 4.000 1515.510 4.280 ;
        RECT 1516.350 4.000 1527.010 4.280 ;
        RECT 1527.850 4.000 1538.050 4.280 ;
        RECT 1538.890 4.000 1549.550 4.280 ;
        RECT 1550.390 4.000 1561.050 4.280 ;
        RECT 1561.890 4.000 1572.550 4.280 ;
        RECT 1573.390 4.000 1584.050 4.280 ;
        RECT 1584.890 4.000 1595.550 4.280 ;
        RECT 1596.390 4.000 1607.050 4.280 ;
        RECT 1607.890 4.000 1618.550 4.280 ;
        RECT 1619.390 4.000 1629.590 4.280 ;
        RECT 1630.430 4.000 1641.090 4.280 ;
        RECT 1641.930 4.000 1652.590 4.280 ;
        RECT 1653.430 4.000 1664.090 4.280 ;
        RECT 1664.930 4.000 1675.590 4.280 ;
        RECT 1676.430 4.000 1687.090 4.280 ;
        RECT 1687.930 4.000 1698.590 4.280 ;
        RECT 1699.430 4.000 1710.090 4.280 ;
        RECT 1710.930 4.000 1721.130 4.280 ;
        RECT 1721.970 4.000 1732.630 4.280 ;
        RECT 1733.470 4.000 1744.130 4.280 ;
        RECT 1744.970 4.000 1755.630 4.280 ;
        RECT 1756.470 4.000 1767.130 4.280 ;
        RECT 1767.970 4.000 1778.630 4.280 ;
        RECT 1779.470 4.000 1790.130 4.280 ;
        RECT 1790.970 4.000 1801.630 4.280 ;
        RECT 1802.470 4.000 1812.670 4.280 ;
        RECT 1813.510 4.000 1824.170 4.280 ;
        RECT 1825.010 4.000 1835.670 4.280 ;
        RECT 1836.510 4.000 1847.170 4.280 ;
        RECT 1848.010 4.000 1858.670 4.280 ;
        RECT 1859.510 4.000 1870.170 4.280 ;
        RECT 1871.010 4.000 1881.670 4.280 ;
        RECT 1882.510 4.000 1893.170 4.280 ;
        RECT 1894.010 4.000 1904.210 4.280 ;
        RECT 1905.050 4.000 1915.710 4.280 ;
        RECT 1916.550 4.000 1927.210 4.280 ;
        RECT 1928.050 4.000 1938.710 4.280 ;
        RECT 1939.550 4.000 1950.210 4.280 ;
        RECT 1951.050 4.000 1961.710 4.280 ;
        RECT 1962.550 4.000 1973.210 4.280 ;
        RECT 1974.050 4.000 1984.710 4.280 ;
        RECT 1985.550 4.000 1995.750 4.280 ;
        RECT 1996.590 4.000 2007.250 4.280 ;
        RECT 2008.090 4.000 2018.750 4.280 ;
        RECT 2019.590 4.000 2030.250 4.280 ;
        RECT 2031.090 4.000 2041.750 4.280 ;
        RECT 2042.590 4.000 2053.250 4.280 ;
        RECT 2054.090 4.000 2064.750 4.280 ;
        RECT 2065.590 4.000 2075.790 4.280 ;
        RECT 2076.630 4.000 2087.290 4.280 ;
        RECT 2088.130 4.000 2098.790 4.280 ;
        RECT 2099.630 4.000 2110.290 4.280 ;
        RECT 2111.130 4.000 2121.790 4.280 ;
        RECT 2122.630 4.000 2133.290 4.280 ;
        RECT 2134.130 4.000 2144.790 4.280 ;
        RECT 2145.630 4.000 2156.290 4.280 ;
        RECT 2157.130 4.000 2167.330 4.280 ;
        RECT 2168.170 4.000 2178.830 4.280 ;
        RECT 2179.670 4.000 2190.330 4.280 ;
        RECT 2191.170 4.000 2201.830 4.280 ;
        RECT 2202.670 4.000 2213.330 4.280 ;
        RECT 2214.170 4.000 2224.830 4.280 ;
        RECT 2225.670 4.000 2236.330 4.280 ;
        RECT 2237.170 4.000 2247.830 4.280 ;
        RECT 2248.670 4.000 2258.870 4.280 ;
        RECT 2259.710 4.000 2270.370 4.280 ;
        RECT 2271.210 4.000 2281.870 4.280 ;
        RECT 2282.710 4.000 2293.370 4.280 ;
        RECT 2294.210 4.000 2304.870 4.280 ;
        RECT 2305.710 4.000 2316.370 4.280 ;
        RECT 2317.210 4.000 2327.870 4.280 ;
        RECT 2328.710 4.000 2339.370 4.280 ;
        RECT 2340.210 4.000 2350.410 4.280 ;
        RECT 2351.250 4.000 2361.910 4.280 ;
        RECT 2362.750 4.000 2373.410 4.280 ;
        RECT 2374.250 4.000 2384.910 4.280 ;
        RECT 2385.750 4.000 2396.410 4.280 ;
        RECT 2397.250 4.000 2407.910 4.280 ;
        RECT 2408.750 4.000 2419.410 4.280 ;
        RECT 2420.250 4.000 2430.910 4.280 ;
        RECT 2431.750 4.000 2441.950 4.280 ;
        RECT 2442.790 4.000 2453.450 4.280 ;
        RECT 2454.290 4.000 2464.950 4.280 ;
        RECT 2465.790 4.000 2476.450 4.280 ;
        RECT 2477.290 4.000 2487.950 4.280 ;
        RECT 2488.790 4.000 2499.450 4.280 ;
        RECT 2500.290 4.000 2510.950 4.280 ;
        RECT 2511.790 4.000 2522.450 4.280 ;
        RECT 2523.290 4.000 2533.490 4.280 ;
        RECT 2534.330 4.000 2544.990 4.280 ;
        RECT 2545.830 4.000 2556.490 4.280 ;
        RECT 2557.330 4.000 2567.990 4.280 ;
        RECT 2568.830 4.000 2579.490 4.280 ;
        RECT 2580.330 4.000 2590.990 4.280 ;
        RECT 2591.830 4.000 2602.490 4.280 ;
        RECT 2603.330 4.000 2613.990 4.280 ;
        RECT 2614.830 4.000 2625.030 4.280 ;
        RECT 2625.870 4.000 2636.530 4.280 ;
        RECT 2637.370 4.000 2648.030 4.280 ;
        RECT 2648.870 4.000 2659.530 4.280 ;
        RECT 2660.370 4.000 2671.030 4.280 ;
        RECT 2671.870 4.000 2682.530 4.280 ;
        RECT 2683.370 4.000 2694.030 4.280 ;
        RECT 2694.870 4.000 2697.800 4.280 ;
      LAYER met3 ;
        RECT 4.000 3247.360 2696.000 3288.645 ;
        RECT 4.000 3245.960 2695.600 3247.360 ;
        RECT 4.000 3140.600 2696.000 3245.960 ;
        RECT 4.000 3139.200 2695.600 3140.600 ;
        RECT 4.000 3034.520 2696.000 3139.200 ;
        RECT 4.000 3033.120 2695.600 3034.520 ;
        RECT 4.000 2927.760 2696.000 3033.120 ;
        RECT 4.000 2926.360 2695.600 2927.760 ;
        RECT 4.000 2821.680 2696.000 2926.360 ;
        RECT 4.000 2820.280 2695.600 2821.680 ;
        RECT 4.000 2714.920 2696.000 2820.280 ;
        RECT 4.000 2713.520 2695.600 2714.920 ;
        RECT 4.000 2608.840 2696.000 2713.520 ;
        RECT 4.000 2607.440 2695.600 2608.840 ;
        RECT 4.000 2502.080 2696.000 2607.440 ;
        RECT 4.000 2500.680 2695.600 2502.080 ;
        RECT 4.000 2396.000 2696.000 2500.680 ;
        RECT 4.000 2394.600 2695.600 2396.000 ;
        RECT 4.000 2289.240 2696.000 2394.600 ;
        RECT 4.000 2287.840 2695.600 2289.240 ;
        RECT 4.000 2182.480 2696.000 2287.840 ;
        RECT 4.000 2181.080 2695.600 2182.480 ;
        RECT 4.000 2076.400 2696.000 2181.080 ;
        RECT 4.000 2075.000 2695.600 2076.400 ;
        RECT 4.000 1969.640 2696.000 2075.000 ;
        RECT 4.000 1968.240 2695.600 1969.640 ;
        RECT 4.000 1863.560 2696.000 1968.240 ;
        RECT 4.000 1862.160 2695.600 1863.560 ;
        RECT 4.000 1756.800 2696.000 1862.160 ;
        RECT 4.000 1755.400 2695.600 1756.800 ;
        RECT 4.000 1650.720 2696.000 1755.400 ;
        RECT 4.400 1649.320 2695.600 1650.720 ;
        RECT 4.000 1543.960 2696.000 1649.320 ;
        RECT 4.000 1542.560 2695.600 1543.960 ;
        RECT 4.000 1437.880 2696.000 1542.560 ;
        RECT 4.000 1436.480 2695.600 1437.880 ;
        RECT 4.000 1331.120 2696.000 1436.480 ;
        RECT 4.000 1329.720 2695.600 1331.120 ;
        RECT 4.000 1225.040 2696.000 1329.720 ;
        RECT 4.000 1223.640 2695.600 1225.040 ;
        RECT 4.000 1118.280 2696.000 1223.640 ;
        RECT 4.000 1116.880 2695.600 1118.280 ;
        RECT 4.000 1011.520 2696.000 1116.880 ;
        RECT 4.000 1010.120 2695.600 1011.520 ;
        RECT 4.000 905.440 2696.000 1010.120 ;
        RECT 4.000 904.040 2695.600 905.440 ;
        RECT 4.000 798.680 2696.000 904.040 ;
        RECT 4.000 797.280 2695.600 798.680 ;
        RECT 4.000 692.600 2696.000 797.280 ;
        RECT 4.000 691.200 2695.600 692.600 ;
        RECT 4.000 585.840 2696.000 691.200 ;
        RECT 4.000 584.440 2695.600 585.840 ;
        RECT 4.000 479.760 2696.000 584.440 ;
        RECT 4.000 478.360 2695.600 479.760 ;
        RECT 4.000 373.000 2696.000 478.360 ;
        RECT 4.000 371.600 2695.600 373.000 ;
        RECT 4.000 266.920 2696.000 371.600 ;
        RECT 4.000 265.520 2695.600 266.920 ;
        RECT 4.000 160.160 2696.000 265.520 ;
        RECT 4.000 158.760 2695.600 160.160 ;
        RECT 4.000 54.080 2696.000 158.760 ;
        RECT 4.000 52.680 2695.600 54.080 ;
        RECT 4.000 9.015 2696.000 52.680 ;
      LAYER met4 ;
        RECT 454.775 17.175 481.440 3167.265 ;
        RECT 483.840 17.175 484.740 3167.265 ;
        RECT 487.140 17.175 558.240 3167.265 ;
        RECT 560.640 17.175 561.540 3167.265 ;
        RECT 563.940 17.175 635.040 3167.265 ;
        RECT 637.440 17.175 638.340 3167.265 ;
        RECT 640.740 17.175 711.840 3167.265 ;
        RECT 714.240 17.175 715.140 3167.265 ;
        RECT 717.540 17.175 788.640 3167.265 ;
        RECT 791.040 17.175 791.940 3167.265 ;
        RECT 794.340 17.175 865.440 3167.265 ;
        RECT 867.840 17.175 868.740 3167.265 ;
        RECT 871.140 17.175 942.240 3167.265 ;
        RECT 944.640 17.175 945.540 3167.265 ;
        RECT 947.940 17.175 1019.040 3167.265 ;
        RECT 1021.440 17.175 1022.340 3167.265 ;
        RECT 1024.740 17.175 1095.840 3167.265 ;
        RECT 1098.240 17.175 1099.140 3167.265 ;
        RECT 1101.540 17.175 1172.640 3167.265 ;
        RECT 1175.040 17.175 1175.940 3167.265 ;
        RECT 1178.340 17.175 1249.440 3167.265 ;
        RECT 1251.840 17.175 1252.740 3167.265 ;
        RECT 1255.140 17.175 1326.240 3167.265 ;
        RECT 1328.640 17.175 1329.540 3167.265 ;
        RECT 1331.940 17.175 1403.040 3167.265 ;
        RECT 1405.440 17.175 1406.340 3167.265 ;
        RECT 1408.740 17.175 1479.840 3167.265 ;
        RECT 1482.240 17.175 1483.140 3167.265 ;
        RECT 1485.540 17.175 1556.640 3167.265 ;
        RECT 1559.040 17.175 1559.940 3167.265 ;
        RECT 1562.340 17.175 1633.440 3167.265 ;
        RECT 1635.840 17.175 1636.740 3167.265 ;
        RECT 1639.140 17.175 1710.240 3167.265 ;
        RECT 1712.640 17.175 1713.540 3167.265 ;
        RECT 1715.940 17.175 1787.040 3167.265 ;
        RECT 1789.440 17.175 1790.340 3167.265 ;
        RECT 1792.740 17.175 1863.840 3167.265 ;
        RECT 1866.240 17.175 1867.140 3167.265 ;
        RECT 1869.540 17.175 1940.640 3167.265 ;
        RECT 1943.040 17.175 1943.940 3167.265 ;
        RECT 1946.340 3159.110 2017.440 3167.265 ;
        RECT 2019.840 3159.350 2020.740 3167.265 ;
        RECT 2023.140 3159.350 2094.240 3167.265 ;
        RECT 2019.840 3159.110 2094.240 3159.350 ;
        RECT 2096.640 3159.350 2097.540 3167.265 ;
        RECT 2099.940 3159.350 2171.040 3167.265 ;
        RECT 2096.640 3159.110 2171.040 3159.350 ;
        RECT 2173.440 3159.350 2174.340 3167.265 ;
        RECT 2176.740 3159.350 2247.840 3167.265 ;
        RECT 2173.440 3159.110 2247.840 3159.350 ;
        RECT 2250.240 3159.350 2251.140 3167.265 ;
        RECT 2253.540 3159.350 2324.640 3167.265 ;
        RECT 2250.240 3159.110 2324.640 3159.350 ;
        RECT 2327.040 3159.350 2327.940 3167.265 ;
        RECT 2330.340 3159.350 2401.440 3167.265 ;
        RECT 2327.040 3159.110 2401.440 3159.350 ;
        RECT 2403.840 3159.350 2404.740 3167.265 ;
        RECT 2407.140 3159.350 2478.240 3167.265 ;
        RECT 2403.840 3159.110 2478.240 3159.350 ;
        RECT 2480.640 3159.350 2481.540 3167.265 ;
        RECT 2483.940 3159.350 2555.040 3167.265 ;
        RECT 2480.640 3159.110 2555.040 3159.350 ;
        RECT 2557.440 3159.350 2558.340 3167.265 ;
        RECT 2560.740 3159.350 2631.840 3167.265 ;
        RECT 2557.440 3159.110 2631.840 3159.350 ;
        RECT 2634.240 3159.350 2635.140 3167.265 ;
        RECT 2637.540 3159.350 2687.945 3167.265 ;
        RECT 2634.240 3159.110 2687.945 3159.350 ;
        RECT 1946.340 2738.810 2687.945 3159.110 ;
        RECT 1946.340 2645.970 2017.440 2738.810 ;
        RECT 2019.840 2738.570 2094.240 2738.810 ;
        RECT 2019.840 2646.210 2020.740 2738.570 ;
        RECT 2023.140 2646.210 2094.240 2738.570 ;
        RECT 2019.840 2645.970 2094.240 2646.210 ;
        RECT 2096.640 2738.570 2171.040 2738.810 ;
        RECT 2096.640 2646.210 2097.540 2738.570 ;
        RECT 2099.940 2646.210 2171.040 2738.570 ;
        RECT 2096.640 2645.970 2171.040 2646.210 ;
        RECT 2173.440 2738.570 2247.840 2738.810 ;
        RECT 2173.440 2646.210 2174.340 2738.570 ;
        RECT 2176.740 2646.210 2247.840 2738.570 ;
        RECT 2173.440 2645.970 2247.840 2646.210 ;
        RECT 2250.240 2738.570 2324.640 2738.810 ;
        RECT 2250.240 2646.210 2251.140 2738.570 ;
        RECT 2253.540 2646.210 2324.640 2738.570 ;
        RECT 2250.240 2645.970 2324.640 2646.210 ;
        RECT 2327.040 2738.570 2401.440 2738.810 ;
        RECT 2327.040 2646.210 2327.940 2738.570 ;
        RECT 2330.340 2646.210 2401.440 2738.570 ;
        RECT 2327.040 2645.970 2401.440 2646.210 ;
        RECT 2403.840 2738.570 2478.240 2738.810 ;
        RECT 2403.840 2646.210 2404.740 2738.570 ;
        RECT 2407.140 2646.210 2478.240 2738.570 ;
        RECT 2403.840 2645.970 2478.240 2646.210 ;
        RECT 2480.640 2738.570 2555.040 2738.810 ;
        RECT 2480.640 2646.210 2481.540 2738.570 ;
        RECT 2483.940 2646.210 2555.040 2738.570 ;
        RECT 2480.640 2645.970 2555.040 2646.210 ;
        RECT 2557.440 2738.570 2631.840 2738.810 ;
        RECT 2557.440 2646.210 2558.340 2738.570 ;
        RECT 2560.740 2646.210 2631.840 2738.570 ;
        RECT 2557.440 2645.970 2631.840 2646.210 ;
        RECT 2634.240 2738.570 2687.945 2738.810 ;
        RECT 2634.240 2646.210 2635.140 2738.570 ;
        RECT 2637.540 2646.210 2687.945 2738.570 ;
        RECT 2634.240 2645.970 2687.945 2646.210 ;
        RECT 1946.340 2225.670 2687.945 2645.970 ;
        RECT 1946.340 2132.830 2017.440 2225.670 ;
        RECT 2019.840 2225.430 2094.240 2225.670 ;
        RECT 2019.840 2133.070 2020.740 2225.430 ;
        RECT 2023.140 2133.070 2094.240 2225.430 ;
        RECT 2019.840 2132.830 2094.240 2133.070 ;
        RECT 2096.640 2225.430 2171.040 2225.670 ;
        RECT 2096.640 2133.070 2097.540 2225.430 ;
        RECT 2099.940 2133.070 2171.040 2225.430 ;
        RECT 2096.640 2132.830 2171.040 2133.070 ;
        RECT 2173.440 2225.430 2247.840 2225.670 ;
        RECT 2173.440 2133.070 2174.340 2225.430 ;
        RECT 2176.740 2133.070 2247.840 2225.430 ;
        RECT 2173.440 2132.830 2247.840 2133.070 ;
        RECT 2250.240 2225.430 2324.640 2225.670 ;
        RECT 2250.240 2133.070 2251.140 2225.430 ;
        RECT 2253.540 2133.070 2324.640 2225.430 ;
        RECT 2250.240 2132.830 2324.640 2133.070 ;
        RECT 2327.040 2225.430 2401.440 2225.670 ;
        RECT 2327.040 2133.070 2327.940 2225.430 ;
        RECT 2330.340 2133.070 2401.440 2225.430 ;
        RECT 2327.040 2132.830 2401.440 2133.070 ;
        RECT 2403.840 2225.430 2478.240 2225.670 ;
        RECT 2403.840 2133.070 2404.740 2225.430 ;
        RECT 2407.140 2133.070 2478.240 2225.430 ;
        RECT 2403.840 2132.830 2478.240 2133.070 ;
        RECT 2480.640 2225.430 2555.040 2225.670 ;
        RECT 2480.640 2133.070 2481.540 2225.430 ;
        RECT 2483.940 2133.070 2555.040 2225.430 ;
        RECT 2480.640 2132.830 2555.040 2133.070 ;
        RECT 2557.440 2225.430 2631.840 2225.670 ;
        RECT 2557.440 2133.070 2558.340 2225.430 ;
        RECT 2560.740 2133.070 2631.840 2225.430 ;
        RECT 2557.440 2132.830 2631.840 2133.070 ;
        RECT 2634.240 2225.430 2687.945 2225.670 ;
        RECT 2634.240 2133.070 2635.140 2225.430 ;
        RECT 2637.540 2133.070 2687.945 2225.430 ;
        RECT 2634.240 2132.830 2687.945 2133.070 ;
        RECT 1946.340 1712.530 2687.945 2132.830 ;
        RECT 1946.340 1619.690 2017.440 1712.530 ;
        RECT 2019.840 1712.290 2094.240 1712.530 ;
        RECT 2019.840 1619.930 2020.740 1712.290 ;
        RECT 2023.140 1619.930 2094.240 1712.290 ;
        RECT 2019.840 1619.690 2094.240 1619.930 ;
        RECT 2096.640 1712.290 2171.040 1712.530 ;
        RECT 2096.640 1619.930 2097.540 1712.290 ;
        RECT 2099.940 1619.930 2171.040 1712.290 ;
        RECT 2096.640 1619.690 2171.040 1619.930 ;
        RECT 2173.440 1712.290 2247.840 1712.530 ;
        RECT 2173.440 1619.930 2174.340 1712.290 ;
        RECT 2176.740 1619.930 2247.840 1712.290 ;
        RECT 2173.440 1619.690 2247.840 1619.930 ;
        RECT 2250.240 1712.290 2324.640 1712.530 ;
        RECT 2250.240 1619.930 2251.140 1712.290 ;
        RECT 2253.540 1619.930 2324.640 1712.290 ;
        RECT 2250.240 1619.690 2324.640 1619.930 ;
        RECT 2327.040 1712.290 2401.440 1712.530 ;
        RECT 2327.040 1619.930 2327.940 1712.290 ;
        RECT 2330.340 1619.930 2401.440 1712.290 ;
        RECT 2327.040 1619.690 2401.440 1619.930 ;
        RECT 2403.840 1712.290 2478.240 1712.530 ;
        RECT 2403.840 1619.930 2404.740 1712.290 ;
        RECT 2407.140 1619.930 2478.240 1712.290 ;
        RECT 2403.840 1619.690 2478.240 1619.930 ;
        RECT 2480.640 1712.290 2555.040 1712.530 ;
        RECT 2480.640 1619.930 2481.540 1712.290 ;
        RECT 2483.940 1619.930 2555.040 1712.290 ;
        RECT 2480.640 1619.690 2555.040 1619.930 ;
        RECT 2557.440 1712.290 2631.840 1712.530 ;
        RECT 2557.440 1619.930 2558.340 1712.290 ;
        RECT 2560.740 1619.930 2631.840 1712.290 ;
        RECT 2557.440 1619.690 2631.840 1619.930 ;
        RECT 2634.240 1712.290 2687.945 1712.530 ;
        RECT 2634.240 1619.930 2635.140 1712.290 ;
        RECT 2637.540 1619.930 2687.945 1712.290 ;
        RECT 2634.240 1619.690 2687.945 1619.930 ;
        RECT 1946.340 1199.390 2687.945 1619.690 ;
        RECT 1946.340 1106.550 2017.440 1199.390 ;
        RECT 2019.840 1199.150 2094.240 1199.390 ;
        RECT 2019.840 1106.790 2020.740 1199.150 ;
        RECT 2023.140 1106.790 2094.240 1199.150 ;
        RECT 2019.840 1106.550 2094.240 1106.790 ;
        RECT 2096.640 1199.150 2171.040 1199.390 ;
        RECT 2096.640 1106.790 2097.540 1199.150 ;
        RECT 2099.940 1106.790 2171.040 1199.150 ;
        RECT 2096.640 1106.550 2171.040 1106.790 ;
        RECT 2173.440 1199.150 2247.840 1199.390 ;
        RECT 2173.440 1106.790 2174.340 1199.150 ;
        RECT 2176.740 1106.790 2247.840 1199.150 ;
        RECT 2173.440 1106.550 2247.840 1106.790 ;
        RECT 2250.240 1199.150 2324.640 1199.390 ;
        RECT 2250.240 1106.790 2251.140 1199.150 ;
        RECT 2253.540 1106.790 2324.640 1199.150 ;
        RECT 2250.240 1106.550 2324.640 1106.790 ;
        RECT 2327.040 1199.150 2401.440 1199.390 ;
        RECT 2327.040 1106.790 2327.940 1199.150 ;
        RECT 2330.340 1106.790 2401.440 1199.150 ;
        RECT 2327.040 1106.550 2401.440 1106.790 ;
        RECT 2403.840 1199.150 2478.240 1199.390 ;
        RECT 2403.840 1106.790 2404.740 1199.150 ;
        RECT 2407.140 1106.790 2478.240 1199.150 ;
        RECT 2403.840 1106.550 2478.240 1106.790 ;
        RECT 2480.640 1199.150 2555.040 1199.390 ;
        RECT 2480.640 1106.790 2481.540 1199.150 ;
        RECT 2483.940 1106.790 2555.040 1199.150 ;
        RECT 2480.640 1106.550 2555.040 1106.790 ;
        RECT 2557.440 1199.150 2631.840 1199.390 ;
        RECT 2557.440 1106.790 2558.340 1199.150 ;
        RECT 2560.740 1106.790 2631.840 1199.150 ;
        RECT 2557.440 1106.550 2631.840 1106.790 ;
        RECT 2634.240 1199.150 2687.945 1199.390 ;
        RECT 2634.240 1106.790 2635.140 1199.150 ;
        RECT 2637.540 1106.790 2687.945 1199.150 ;
        RECT 2634.240 1106.550 2687.945 1106.790 ;
        RECT 1946.340 686.250 2687.945 1106.550 ;
        RECT 1946.340 593.410 2017.440 686.250 ;
        RECT 2019.840 686.010 2094.240 686.250 ;
        RECT 2019.840 593.650 2020.740 686.010 ;
        RECT 2023.140 593.650 2094.240 686.010 ;
        RECT 2019.840 593.410 2094.240 593.650 ;
        RECT 2096.640 686.010 2171.040 686.250 ;
        RECT 2096.640 593.650 2097.540 686.010 ;
        RECT 2099.940 593.650 2171.040 686.010 ;
        RECT 2096.640 593.410 2171.040 593.650 ;
        RECT 2173.440 686.010 2247.840 686.250 ;
        RECT 2173.440 593.650 2174.340 686.010 ;
        RECT 2176.740 593.650 2247.840 686.010 ;
        RECT 2173.440 593.410 2247.840 593.650 ;
        RECT 2250.240 686.010 2324.640 686.250 ;
        RECT 2250.240 593.650 2251.140 686.010 ;
        RECT 2253.540 593.650 2324.640 686.010 ;
        RECT 2250.240 593.410 2324.640 593.650 ;
        RECT 2327.040 686.010 2401.440 686.250 ;
        RECT 2327.040 593.650 2327.940 686.010 ;
        RECT 2330.340 593.650 2401.440 686.010 ;
        RECT 2327.040 593.410 2401.440 593.650 ;
        RECT 2403.840 686.010 2478.240 686.250 ;
        RECT 2403.840 593.650 2404.740 686.010 ;
        RECT 2407.140 593.650 2478.240 686.010 ;
        RECT 2403.840 593.410 2478.240 593.650 ;
        RECT 2480.640 686.010 2555.040 686.250 ;
        RECT 2480.640 593.650 2481.540 686.010 ;
        RECT 2483.940 593.650 2555.040 686.010 ;
        RECT 2480.640 593.410 2555.040 593.650 ;
        RECT 2557.440 686.010 2631.840 686.250 ;
        RECT 2557.440 593.650 2558.340 686.010 ;
        RECT 2560.740 593.650 2631.840 686.010 ;
        RECT 2557.440 593.410 2631.840 593.650 ;
        RECT 2634.240 686.010 2687.945 686.250 ;
        RECT 2634.240 593.650 2635.140 686.010 ;
        RECT 2637.540 593.650 2687.945 686.010 ;
        RECT 2634.240 593.410 2687.945 593.650 ;
        RECT 1946.340 173.110 2687.945 593.410 ;
        RECT 1946.340 17.175 2017.440 173.110 ;
        RECT 2019.840 172.870 2094.240 173.110 ;
        RECT 2019.840 17.175 2020.740 172.870 ;
        RECT 2023.140 17.175 2094.240 172.870 ;
        RECT 2096.640 172.870 2171.040 173.110 ;
        RECT 2096.640 17.175 2097.540 172.870 ;
        RECT 2099.940 17.175 2171.040 172.870 ;
        RECT 2173.440 172.870 2247.840 173.110 ;
        RECT 2173.440 17.175 2174.340 172.870 ;
        RECT 2176.740 17.175 2247.840 172.870 ;
        RECT 2250.240 172.870 2324.640 173.110 ;
        RECT 2250.240 17.175 2251.140 172.870 ;
        RECT 2253.540 17.175 2324.640 172.870 ;
        RECT 2327.040 172.870 2401.440 173.110 ;
        RECT 2327.040 17.175 2327.940 172.870 ;
        RECT 2330.340 17.175 2401.440 172.870 ;
        RECT 2403.840 172.870 2478.240 173.110 ;
        RECT 2403.840 17.175 2404.740 172.870 ;
        RECT 2407.140 17.175 2478.240 172.870 ;
        RECT 2480.640 172.870 2555.040 173.110 ;
        RECT 2480.640 17.175 2481.540 172.870 ;
        RECT 2483.940 17.175 2555.040 172.870 ;
        RECT 2557.440 172.870 2631.840 173.110 ;
        RECT 2557.440 17.175 2558.340 172.870 ;
        RECT 2560.740 17.175 2631.840 172.870 ;
        RECT 2634.240 172.870 2687.945 173.110 ;
        RECT 2634.240 17.175 2635.140 172.870 ;
        RECT 2637.540 17.175 2687.945 172.870 ;
  END
END top_level_bASIC
END LIBRARY

